Mirinae �                �0! <  �.!     �K  p   p                                              ������                                                                                                                                                                                                                                                                                                                                                                                                                      T T i W W B W5 B2 W B W6 D3 B2 W s B W4 W5 D i W W i i2 i i        ��   	 2                    �  X    $                     �zb���� � ������������               ��  	  2                 
     $    #                    �zb���� � ������������               �� 	   2    #                0  `    !                    �zb���� � ������������               ��	    2    (                N  �                        �zb���� � ������������               ��    2    -                l  �                       �zb���� � ������������               ��    2    2                �                         �zb���� � ������������               ��    2    7                �  P                       �zb���� � ������������               ��    2    <                �  �                       �zb���� � ������������               ��    2    A                �  �                       �zb���� � ������������               ��    2    F                          	               �zb���� � ������������               ��    2    4 #              z  n
    "                   ������� � ������������              ��    2    9 '              �  "    !                  ������� � ������������              ��   ! 2    > +              �  �                      ������� � ������������              �� ! " % 2    C /               .  �                     ������� � ������������              �� % & ) 2    H 3           !   j  >                     ������� � ������������              ��! ) * - 2    M 7           #   �  �                     ������� � ������������              ��$ - . 1 2    R ;           %   �  �                     ������� � ������������              ��' 1 2 5 2    W ?           '     Z                     ������� � ������������              ��* 5 6 9 2    \ C           )   Z                       ������� � ������������              ��- 9 : = 2    a G           *   �  �        	             ������� � ������������              ��% 3 3 7 2    N 4          B   �                          b������ � ������������              ��* 8 8 = 2    S 8 !         F   �  �                      b������ � ������������              ��/ = = C 2    X < $         J   :  �                      b������ � ������������              ��4 B B I 2    ] @ '         M   �  P                     b������ � ������������              ��9 G G O 2    b D *         Q   �  �                     b������ � ������������              ��> L L U 2    g H -         T   H   !                     b������ � ������������              ��C Q Q [ 2    l L 0         X   �  �"                     b������ � ������������              ��H V V a 2    q P 3         \   �  �#                     b������ � ������������              ��M [ [ g 2    v T 6         _   V	  X%                     b������ � ������������              ��R ` ` m 2    { X 9         c   �	  �&        	             b������ � ������������              ��F V T d 2    g D &        �     x7                       �q����� � ������������              ��L ] [ k 2    l H )        �   �  �9                      �q����� � ������������              ��R d b r 2    q L ,         �     (<                      �q����� � ������������              ��X k i y 2    v P / #       �   �  �>                     �q����� � ������������              ��^ r p � 2    { T 2 &       �   �  �@                     �q����� � ������������              ��d y w � 2    � X 5 )       �   p  0C                     �q����� � ������������              ��j � ~ � 2    � \ 8 ,       �   �  �E                     �q����� � ������������              ��p � � � 2    � ` ; /       �   `  �G                     �q����� � ������������              ��v � � � 2    � d > 2       �   �  8J                     �q����� � ������������              ��| � � � 2    � h A 5       �   P  �L        	             �q����� � ������������              ��k � � � 2     S - !         0   g                       ֚c���� � ������������              ��s � � � 2    � W 0 $         �  �j                      ֚c���� � ������������              ��{ � � � 2    � [ 3 '         \  (n                      ֚c���� � ������������              ��� � � � 2    � _ 6 *       #  �  �q                     ֚c���� � ������������              ��� � � � 2    � c 9 -       ,  �  0u                     ֚c���� � ������������              ��� � � � 2    � g < 0       5    �x                     ֚c���� � ������������              ��� � � � 2    � k ? 3       >  �  8|                     ֚c���� � ������������              ��� � � � 2    � o B 6       G  J  �                     ֚c���� � ������������              ��� � � � 2    � s E 9       P  �  @�                     ֚c���� � ������������              ��� � � � 2    � w H <       Y  v  Ć        	             ֚c���� � ������������              ��� � � � 2    � b 4 (       �  �  ��                       ~S����� � ������������              ��� � � � 2    � g 7 +       �  �  ��                      ~S����� � ������������              ��� � � � 2    � l : .       �  6  z�                      ~S����� � ������������              ��� � � � 2    � q = 1       �  �  f�                     ~S����� � ������������              ��� � � 2    � v @ 4       �  �  R�                     ~S����� � ������������              ��� � � 2    � { C 7       �  R  >�                     ~S����� � ������������              ��� � � 2    � � F :           *�                     ~S����� � ������������              ��� � � "2    � � I =         �  �                     ~S����� � ������������              ��� -2    � � L @       !  n  �                     ~S����� � ������������              ��� 82    � � O C       -  "  ��        	             ~S����� � ������������              ��� � � #2    � z : .       �  �!  �                      BE����� � �����  �                ��� /2    �  > 2       �  �"                        BE����� � �����  �                ��� ;2    � � B 6       �  �#  �                     BE����� � �����  �                ��� G2    � � F :       �  h$  @#                    BE����� � �����  �                ��� #)S2    � � J >       �  :%  �)                    BE����� � �����  �                ��	.5_2    � � N B         &  `0                    BE����� � �����  �                ��9Ak2    � � R F         �&  �6                    BE����� � �����  �                ��DMw2    � � V J       ,  �'  �=                    BE����� � �����  �                ��'OY�2    � � Z N       =  �(  D                    BE����� � �����  �                ��1Ze�2    � � ^ R       N  T)  �J       	             BE����� � �����  �                ��	    2    (                �  H    $                  ������� � ������������              ��    2    -                      #                 ������� � ������������              ��    2    2                   @    !                 ������� � ������������              ��   	 2    7                >  |                     ������� � ������������              ��  	  2    <                \  �                    ������� � ������������              ��    2    A                z  �                    ������� � ������������              ��    2    F                �  0                    ������� � ������������              ��    2    K                �  l                    ������� � ������������              ��    2    P                �  �                    ������� � ������������              ��    2    U                �  �        	            ������� � ������������              ��    2    C 2           !   j  >    "                  ������� � ������������              ��    2    H 6           #   �  �    !                 ������� � ������������              ��  #   2    M :           %   �  �                     ������� � ������������              ��$ '   2    R >           '     Z                    ������� � ������������              ��( +   2    W B           )   Z                      ������� � ������������              ��, /  " 2    \ F           *   �  �                    ������� � ������������              ��0 3 " % 2    a J           ,   �  v                    ������� � ������������              ��4 7 % ( 2    f N           .     *                    ������� � ������������              ��8 ; ( + 2    k R           0   J  �                    ������� � ������������              ��< ? + . 2    p V           2   �  �        	            ������� � ������������              ��5 9 # ' 2    ] C          L   v  �                  	     ������� � ������������	              ��; ? ' , 2    b G !         P   �  @                	     ������� � ������������	              ��A E + 1 2    g K $         S   *  �                 	     ������� � ������������	              ��G K / 6 2    l O '         W   �  "                	    ������� � ������������	              ��M Q 3 ; 2    q S *         Z   �  x#                	    ������� � ������������	              ��S W 7 @ 2    v W -         ^   8	  �$                	    ������� � ������������	              ��Y ] ; E 2    { [ 0         b   �	  H&                	    ������� � ������������	              ��_ c ? J 2    � _ 3         e   �	  �'                	    ������� � ������������	              ��e i C O 2    � c 6         i   F
  )                	    ������� � ������������	              ��k o G T 2    � g 9         l   �
  �*        	        	    ������� � ������������	              ��` f : J 2    v S &        �     (<                 
     ��@���� � ������������
              ��g n @ P 2    { W )        �   �  �>                
     ��@���� � ������������
              ��n v F V 2    � [ ,         �   �  �@                
     ��@���� � ������������
              ��u ~ L \ 2    � _ / #       �   p  0C                
    ��@���� � ������������
              ��| � R b 2    � c 2 &       �   �  �E                
    ��@���� � ������������
              ��� � X h 2    � g 5 )       �   `  �G                
    ��@���� � ������������
              ��� � ^ n 2    � k 8 ,       �   �  8J                
    ��@���� � ������������
              ��� � d t 2    � o ; /       �   P  �L                
    ��@���� � ������������
              ��� � j z 2    � s > 2       �   �  �N                
    ��@���� � ������������
              ��� � p � 2    � w A 5       �   @  @Q        	        
    ��@���� � ������������
              ��� � _ q 2    � b - !            �l                      ������� � ������������              ��� � f y 2    � f 0 $         �  Dp                     ������� � ������������              ��� � m � 2    � j 3 '       (  L  �s                     ������� � ������������              ��� � t � 2    � n 6 *       1  �  Lw                    ������� � ������������              ��� � { � 2    � r 9 -       :  x  �z                    ������� � ������������              ��� � � � 2    � v < 0       C    T~                    ������� � ������������              ��� � � � 2    � z ? 3       L  �  ؁                    ������� � ������������              ��� � � � 2    � ~ B 6       U  :  \�                    ������� � ������������              ��� � � � 2    � � E 9       ^  �  ��                    ������� � ������������              ��� � � � 2    � � H <       g  f  d�        	            ������� � ������������              ��� � � � 2    � q 4 (       �  �  2�                      k������ � ������������              ��� � � � 2    � v 7 +       �  r  �                     k������ � ������������              ��� � � � 2    � { : .       �  &  
�                     k������ � ������������              ��� � � 2    � � = 1       �  �  ��                    k������ � ������������              ��� � � 2    � � @ 4       �  �  ��                    k������ � ������������              ��� � 2    � � C 7         B  ��                    k������ � ������������              ��#� � 2    � � F :         �  ��                    k������ � ������������              ��.� � 2    � � I =       %  �  ��                    k������ � ������������              ��%9� � 2    � � L @       2  ^  ��                    k������ � ������������              ��0D� � 2    � � O C       >     ~�        	            k������ � ������������              ��/� � 2    � � : .       �  �"                       ������� � �����  �                ��%<� � 2    � � > 2       �  �#  �                    ������� � �����  �                ��1I� � 2    � � B 6       �  �$  0$                    ������� � �����  �                ��=V� � 2    � � F :       �  X%  �*                   ������� � �����  �                ��Ic� 	2    � � J >         *&  P1                   ������� � �����  �                ��Up� 2    � � N B         �&  �7                   ������� � �����  �                ��a}� 2    � � R F       /  �'  p>                   ������� � �����  �                ��m�� '2    � � V J       @  �(   E                   ������� � �����  �                ��y�12    � Z N       P  r)  �K                   ������� � �����  �                ����;2    � ^ R       a  D*   R       	            ������� � �����  �                ��    2                   0  �    $   ,       *        ��{���� � ������������              �� 	  	 2    "   "            N  �    #   ,      *        ��{���� � ������������              ��	  	  2    &   &            l  �    !   ,      *        ��{���� � ������������              ��    2    *   *            �          ,      *       ��{���� � ������������              ��    2    .   .            �  P       ,      *       ��{���� � ������������              ��    2    2   2            �  �       ,      *       ��{���� � ������������              ��    2    6   6            �  �       ,      *       ��{���� � ������������              ��    2    :   :                     ,      *       ��{���� � ������������              ��    2    >   >               @       ,      *       ��{���� � ������������              ��    2    B   B            >  |       , 	     *       ��{���� � ������������              ��    2    / ( /            �  "    "   -       +        ������� � ������������              ��    2    3 * 3            �  �    !   -      +        ������� � ������������              ��    2    7 , 7             .  �       -      +        ������� � ������������              �� #  # 2    ; . ;         !   j  >       -      +       ������� � ������������              ��  '   ' 2    ? 0 ?         #   �  �       -      +       ������� � ������������              ��# + # + 2    C 2 C         %   �  �       -      +       ������� � ������������              ��& / & / 2    G 4 G         '     Z       -      +       ������� � ������������              ��) 3 ) 3 2    K 6 K         )   Z         -      +       ������� � ������������              ��, 7 , 7 2    O 8 O         *   �  �       -      +       ������� � ������������              ��/ ; / ; 2    S : S         ,   �  v       - 	     +       ������� � ������������              ��' 5 ' 5 2    @ & @        E   �          .       ,        ������� � ������������              ��, : , : 2    E ) E        H     p       .      ,        ������� � ������������              ��1 ? 1 ? 2    J , J         L   v  �       .      ,        ������� � ������������              ��6 D 6 D 2    O / O #       P   �  @       .      ,       ������� � ������������              ��; I ; I 2    T 2 T &       S   *  �        .      ,       ������� � ������������              ��@ N @ N 2    Y 5 Y )       W   �  "       .      ,       ������� � ������������              ��E S E S 2    ^ 8 ^ ,       Z   �  x#       .      ,       ������� � ������������              ��J X J X 2    c ; c /       ^   8	  �$       .      ,       ������� � ������������              ��O ] O ] 2    h > h 2       b   �	  H&       .      ,       ������� � ������������              ��T b T b 2    m A m 5       e   �	  �'       . 	     ,       ������� � ������������              ��H X H X 2    Z . Z "       �   T  �8       /       -        ������� � ������������              ��N _ N _ 2    _ 1 _ %       �   �  �:       /      -        ������� � ������������              ��T f T f 2    d 4 d (       �   D  T=       /      -        ������� � ������������              ��Z m Z m 2    i 7 i +       �   �  �?       /      -       ������� � ������������              ��` t ` t 2    n : n .       �   4  B       /      -       ������� � ������������              ��f { f { 2    s = s 1       �   �  \D       /      -       ������� � ������������              ��l � l � 2    x @ x 4       �   $  �F       /      -       ������� � ������������              ��r � r � 2    } C } 7       �   �  I       /      -       ������� � ������������              ��x � x � 2    � F � :       �     dK       /      -       ������� � ������������              ��~ � ~ � 2    � I � =       �   �  �M       / 	     -       ������� � ������������              ��m � m � 2    s 5 s )         l  �h       0       .        D�n���� � ������������              ��u � u � 2    x 8 x ,           l       0      .        D�n���� � ������������              ��} � } � 2    } ; } /         �  �o       0      .        D�n���� � ������������              ��� � � � 2    � > � 2       &  .  s       0      .       D�n���� � ������������              ��� � � � 2    � A � 5       /  �  �v       0      .       D�n���� � ������������              ��� � � � 2    � D � 8       8  Z  z       0      .       D�n���� � ������������              ��� � � � 2    � G � ;       A  �  �}       0      .       D�n���� � ������������              ��� � � � 2    � J � >       J  �  $�       0      .       D�n���� � ������������              ��� � � � 2    � M � A       S    ��       0      .       D�n���� � ������������              ��� � � � 2    � P � D       \  �  ,�       0 	     .       D�n���� � ������������              ��� � � � 2    � < � 0       �  
  F�       1       /        ������� � ������������              ��� � � � 2    � ? � 3       �  �  2�       1      /        ������� � ������������              ��� � � � 2    � B � 6       �  r  �       1      /        ������� � ������������              ��� � � � 2    � E � 9       �  &  
�       1      /       ������� � ������������              ��� � � � 2    � H � <       �  �  ��       1      /       ������� � ������������              ��� � � � 2    � K � ?       �  �  ��       1      /       ������� � ������������              ��� � 2    � N � B         B  ��       1      /       ������� � ������������              ��� � 2    � Q � E         �  ��       1      /       ������� � ������������              ��� � 2    � T � H       %  �  ��       1      /       ������� � ������������              ��� #� #2    � W � K       2  ^  ��       1 	     /       ������� � ������������              ��� � 2    � B � 6       �  ."  p      2       0        Ǥ^���� � �����  �                ��� � 2    � F � :       �   #         2      0        Ǥ^���� � �����  �                ��� %� %2    � J � >       �  �#  �      2      0        Ǥ^���� � �����  �                ��112    � N � B       �  �$   %      2      0       Ǥ^���� � �����  �                ��==2    � R � F       �  v%  �+      2      0       Ǥ^���� � �����  �                ��II2    � V � J         H&  @2      2      0       Ǥ^���� � �����  �                ��%U%U2    � Z � N          '  �8      2      0       Ǥ^���� � �����  �                ��0a0a2    � ^ � R       1  �'  `?      2      0       Ǥ^���� � �����  �                ��;m;m2    � b � V       B  �(  �E      2      0       Ǥ^���� � �����  �                ��FyFy2    � f � Z       S  �)  �L      2 	     0       Ǥ^���� � �����  �                �� 	   2    #                �      $   B       ?        u}����� � ������������              ��	    2    (                �  �    #   B      ?        u}����� � ������������              ��   	 2    -                �  �    !   B      ?        u}����� � ������������              ��  	  2    2                          B      ?       u}����� � ������������              ��    2    7                   @       B      ?       u}����� � ������������              ��    2    <                >  |       B      ?       u}����� � ������������              ��    2    A                \  �       B      ?       u}����� � ������������              ��    2    F                z  �       B      ?       u}����� � ������������              ��    2    K                �  0       B      ?       u}����� � ������������              ��    2    P                �  l       B 	     ?       u}����� � ������������              ��    2    > -               .  �    "   C       @        ��w���� � ������������              ��    2    C 1           !   j  >    !   C      @        ��w���� � ������������              �� !   2    H 5           #   �  �       C      @        ��w���� � ������������              ��" %  ! 2    M 9           %   �  �       C      @       ��w���� � ������������              ��& )  % 2    R =           '     Z       C      @       ��w���� � ������������              ��* - ! ) 2    W A           )   Z         C      @       ��w���� � ������������              ��. 1 $ - 2    \ E           *   �  �       C      @       ��w���� � ������������              ��2 5 ' 1 2    a I           ,   �  v       C      @       ��w���� � ������������              ��6 9 * 5 2    f M           .     *       C      @       ��w���� � ������������              ��: = - 9 2    k Q           0   J  �       C 	     @       ��w���� � ������������              ��3 7 % 3 2    X >          J   :  �        D       A        ������� � ������������              ��8 = * 8 2    ] B !         M   �  P       D      A        ������� � ������������              ��= C / = 2    b F $         Q   �  �       D      A        ������� � ������������              ��B I 4 B 2    g J '         T   H   !       D      A       ������� � ������������              ��G O 9 G 2    l N *         X   �  �"       D      A       ������� � ������������              ��L U > L 2    q R -         \   �  �#       D      A       ������� � ������������              ��Q [ C Q 2    v V 0         _   V	  X%       D      A       ������� � ������������              ��V a H V 2    { Z 3         c   �	  �&       D      A       ������� � ������������              ��[ g M [ 2    � ^ 6         f   

  ((       D      A       ������� � ������������              ��` m R ` 2    � b 9         j   d
  �)       D 	     A       ������� � ������������              ��T d F V 2    q N &        �   �  �:       E       B        R������ � ������������              ��[ k L ] 2    v R )        �   D  T=       E      B        R������ � ������������              ��b r R d 2    { V ,         �   �  �?       E      B        R������ � ������������              ��i y X k 2    � Z / #       �   4  B       E      B       R������ � ������������              ��p � ^ r 2    � ^ 2 &       �   �  \D       E      B       R������ � ������������              ��w � d y 2    � b 5 )       �   $  �F       E      B       R������ � ������������              ��~ � j � 2    � f 8 ,       �   �  I       E      B       R������ � ������������              ��� � p � 2    � j ; /       �     dK       E      B       R������ � ������������              ��� � v � 2    � n > 2       �   �  �M       E      B       R������ � ������������              ��� � | � 2    � r A 5       �     P       E 	     B       R������ � ������������              ��� � k � 2    � ] - !         �  Xk       F       C        ������� � ������������              ��� � s � 2    � a 0 $         z  �n       F      C        ������� � ������������              ��� � { � 2    � e 3 '       $    `r       F      C        ������� � ������������              ��� � � � 2    � i 6 *       -  �  �u       F      C       ������� � ������������              ��� � � � 2    � m 9 -       6  <  hy       F      C       ������� � ������������              ��� � � � 2    � q < 0       ?  �  �|       F      C       ������� � ������������              ��� � � � 2    � u ? 3       H  h  p�       F      C       ������� � ������������              ��� � � � 2    � y B 6       Q  �  �       F      C       ������� � ������������              ��� � � � 2    � } E 9       Z  �  x�       F      C       ������� � ������������              ��� � � � 2    � � H <       c  *  ��       F 	     C       ������� � ������������              ��� � � � 2    � l 4 (       �  �  ��       G       D        눮���� � ������������              ��� � � � 2    � q 7 +       �  6  z�       G      D        눮���� � ������������              ��� � � � 2    � v : .       �  �  f�       G      D        눮���� � ������������              ��� � � � 2    � { = 1       �  �  R�       G      D       눮���� � ������������              ��� � � 2    � � @ 4       �  R  >�       G      D       눮���� � ������������              ��� � � 2    � � C 7           *�       G      D       눮���� � ������������              ��� � � 2    � � F :         �  �       G      D       눮���� � ������������              ��� "� � 2    � � I =       !  n  �       G      D       눮���� � ������������              ��-� 2    � � L @       -  "  ��       G      D       눮���� � ������������              ��8� 2    � � O C       :  �  ��       G 	     D       눮���� � ������������              ��� #� � 2    � � : .       �  �"  0      H       E        dc����� � �����  �                ��/� 2    � � > 2       �  x#  �      H      E        dc����� � �����  �                ��;� 2    � � B 6       �  J$  P"      H      E        dc����� � �����  �                ��G� 2    � � F :       �  %  �(      H      E       dc����� � �����  �                ��)S� #2    � � J >         �%  p/      H      E       dc����� � �����  �                ��5_	.2    � � N B         �&   6      H      E       dc����� � �����  �                ��Ak92    � � R F       *  �'  �<      H      E       dc����� � �����  �                ��MwD2    � � V J       ;  d(   C      H      E       dc����� � �����  �                ��Y�'O2    � � Z N       L  6)  �I      H      E       dc����� � �����  �                ��e�1Z2    � ^ R       \  *  @P      H 	     E       dc����� � �����  �                ��  	  2                  �      $   X       T        �y����� � ������������              ��    2      #         	   �  �    #   X      T        �y����� � ������������              ��    2      (         
   �  �    !   X      T        �y����� � ������������              �� 	   2     " -         
     $        X      T       �y����� � ������������              ��	    2     % 2            0  `       X      T       �y����� � ������������              ��    2     ( 7            N  �       X      T       �y����� � ������������              ��    2      + <            l  �       X      T       �y����� � ������������              ��    2    " . A            �         X      T       �y����� � ������������              ��    2    $ 1 F            �  P       X      T       �y����� � ������������              ��    2    & 4 K            �  �       X 	     T       �y����� � ������������              ��    2     ! 9           >  �	    "   Y       U        ZY����� � ������������              ��    2     $ >           z  n
    !   Y      U        ZY����� � ������������              ��    # 2     ' C           �  "       Y      U        ZY����� � ������������              ��  $ ' 2     * H            �  �       Y      U       ZY����� � ������������              ��  ( + 2     - M "           .  �       Y      U       ZY����� � ������������              �� " , / 2    " 0 R $       !   j  >       Y      U       ZY����� � ������������              ��" % 0 3 2    % 3 W &       #   �  �       Y      U       ZY����� � ������������              ��% ( 4 7 2    ( 6 \ (       %   �  �       Y      U       ZY����� � ������������              ��( + 8 ; 2    + 9 a *       '     Z       Y      U       ZY����� � ������������              ��+ . < ? 2    . < f ,       )   Z         Y 	     U       ZY����� � ������������              ��# ' 5 9 2     ( S        @   J  (        Z       V        ��s���� � ������������              ��' , ; ? 2     , X        D   �  �       Z      V        ��s���� � ������������              ��+ 1 A E 2    ! 0 ]        G   �  �       Z      V        ��s���� � ������������              ��/ 6 G K 2    $ 4 b !       K   X  `       Z      V       ��s���� � ������������              ��3 ; M Q 2    ' 8 g $       N   �  �       Z      V       ��s���� � ������������              ��7 @ S W 2    * < l '       R     0        Z      V       ��s���� � ������������              ��; E Y ] 2    - @ q *       V   f  �!       Z      V       ��s���� � ������������              ��? J _ c 2    0 D v -       Y   �   #       Z      V       ��s���� � ������������              ��C O e i 2    3 H { 0       ]   	  h$       Z      V       ��s���� � ������������              ��G T k o 2    6 L � 3       `   t	  �%       Z 	     V       ��s���� � ������������              ��: J ` f 2    # 9 l         �   �
  L6       [       W        �e����� � ������������              ��@ P g n 2    & = q #       �   T  �8       [      W        �e����� � ������������              ��F V n v 2    ) A v &       �   �  �:       [      W        �e����� � ������������              ��L \ u ~ 2    , E { )       �   D  T=       [      W       �e����� � ������������              ��R b | � 2    / I � ,       �   �  �?       [      W       �e����� � ������������              ��X h � � 2    2 M � /       �   4  B       [      W       �e����� � ������������              ��^ n � � 2    5 Q � 2       �   �  \D       [      W       �e����� � ������������              ��d t � � 2    8 U � 5       �   $  �F       [      W       �e����� � ������������              ��j z � � 2    ; Y � 8       �   �  I       [      W       �e����� � ������������              ��p � � � 2    > ] � ;       �     dK       [ 	     W       �e����� � ������������              ��_ q � � 2    * I � '         �  �e       \       X         ������ � ������������               ��f y � � 2    - M � *         �  <i       \      X         ������ � ������������               ��m � � � 2    0 Q � -            �l       \      X         ������ � ������������               ��t � � � 2    3 U � 0         �  Dp       \      X        ������ � ������������               ��{ � � � 2    6 Y � 3       (  L  �s       \      X        ������ � ������������               ��� � � � 2    9 ] � 6       1  �  Lw       \      X        ������ � ������������               ��� � � � 2    < a � 9       :  x  �z       \      X        ������ � ������������               ��� � � � 2    ? e � <       C    T~       \      X        ������ � ������������               ��� � � � 2    B i � ?       L  �  ؁       \      X        ������ � ������������               ��� � � � 2    E m � B       U  :  \�       \ 	     X        ������ � ������������               ��� � � � 2    1 X � .       �  �  ��       ]       Y   !     c������ � ������������!              ��� � � � 2    5 \ � 1       �  F  �       ]      Y   !     c������ � ������������!              ��� � � � 2    9 ` � 4       �  �  ֵ       ]      Y   !     c������ � ������������!              ��� � � 2    = d � 7       �  �  º       ]      Y   !    c������ � ������������!              ��� � � 2    A h � :       �  b  ��       ]      Y   !    c������ � ������������!              ��� � 2    E l � =       �    ��       ]      Y   !    c������ � ������������!              ��� � #2    I p � @         �  ��       ]      Y   !    c������ � ������������!              ��� � .2    M t � C         ~  r�       ]      Y   !    c������ � ������������!              ��� � %92    Q x � F         2  ^�       ]      Y   !    c������ � ������������!              ��� � 0D2    U | � I       )  �  J�       ] 	     Y   !    c������ � ������������!              ��� � /2    A g � 4       �  �!  �      ^       Z   "     ��c���� � �����  �  "              ��� � %<2    E l � 8       �  �"  @      ^      Z   "     ��c���� � �����  �  "              ��� � 1I2    I q � <       �  Z#  �      ^      Z   "     ��c���� � �����  �  "              ��� � =V2    M v � @       �  ,$  `!      ^      Z   "    ��c���� � �����  �  "              ��� 	Ic2    Q { � D       �  �$  �'      ^      Z   "    ��c���� � �����  �  "              ��� Up2    U � � H         �%  �.      ^      Z   "    ��c���� � �����  �  "              ��� a}2    Y � � L         �&  5      ^      Z   "    ��c���� � �����  �  "              ��� 'm�2    ] � � P       (  t'  �;      ^      Z   "    ��c���� � �����  �  "              ��1y�2    a � � T       8  F(  0B      ^      Z   "    ��c���� � �����  �  "              ��;��2    e � � X       I  )  �H      ^ 	     Z   "    ��c���� � �����  �  "                   
2                   l  �    $   r       l   #     ������� � ������������#                   
2        "            �      #   r      l   #     ������� � ������������#                
  
 
2    $   &            �  P    !   r      l   #     ������� � ������������#               
  
  
2    (   *            �  �        r      l   #    ������� � ������������#                   
2    ,   .            �  �       r      l   #    ������� � ������������#                   
2    0   2                     r      l   #    ������� � ������������#                   
2    4   6               @       r      l   #    ������� � ������������#                   
2    8   :            >  |       r      l   #    ������� � ������������#                   
2    <   >            \  �       r      l   #    ������� � ������������#                   
2    @   B            z  �       r 	     l   #    ������� � ������������#                   
2    - ( /            �  �    "   s       m   $     ������� � ������������$                   
2    1 * 3             .  �    !   s      m   $     ������� � ������������$                   
2    5 , 7         !   j  >       s      m   $     ������� � ������������$                "  " 
2    9 . ;         #   �  �       s      m   $    ������� � ������������$                &  & 
2    = 0 ?         %   �  �       s      m   $    ������� � ������������$               " * " * 
2    A 2 C         '     Z       s      m   $    ������� � ������������$               % . % . 
2    E 4 G         )   Z         s      m   $    ������� � ������������$               ( 2 ( 2 
2    I 6 K         *   �  �       s      m   $    ������� � ������������$               + 6 + 6 
2    M 8 O         ,   �  v       s      m   $    ������� � ������������$               . : . : 
2    Q : S         .     *       s 	     m   $    ������� � ������������$               & 4 & 4 
2    > & @        G   �  �        t       n   %     ������� � ������������%               + 9 + 9 
2    C ) E        K   X  `       t      n   %     ������� � ������������%               0 > 0 > 
2    H , J         N   �  �       t      n   %     ������� � ������������%               5 C 5 C 
2    M / O #       R     0        t      n   %    ������� � ������������%               : H : H 
2    R 2 T &       V   f  �!       t      n   %    ������� � ������������%               ? M ? M 
2    W 5 Y )       Y   �   #       t      n   %    ������� � ������������%               D R D R 
2    \ 8 ^ ,       ]   	  h$       t      n   %    ������� � ������������%               I W I W 
2    a ; c /       `   t	  �%       t      n   %    ������� � ������������%               N \ N \ 
2    f > h 2       d   �	  8'       t      n   %    ������� � ������������%               S a S a 
2    k A m 5       h   (
  �(       t 	     n   %    ������� � ������������%               G W G W 
2    X . Z "       �   �  �9       u       o   &     ������� � ������������&               M ^ M ^ 
2    ] 1 _ %       �     (<       u      o   &     ������� � ������������&               S e S e 
2    b 4 d (       �   �  �>       u      o   &     ������� � ������������&               Y l Y l 
2    g 7 i +       �   �  �@       u      o   &    ������� � ������������&               _ s _ s 
2    l : n .       �   p  0C       u      o   &    ������� � ������������&               e z e z 
2    q = s 1       �   �  �E       u      o   &    ������� � ������������&               k � k � 
2    v @ x 4       �   `  �G       u      o   &    ������� � ������������&               q � q � 
2    { C } 7       �   �  8J       u      o   &    ������� � ������������&               w � w � 
2    � F � :       �   P  �L       u      o   &    ������� � ������������&               } � } � 
2    � I � =       �   �  �N       u 	     o   &    ������� � ������������&               l � l � 
2    q 5 s )         �  �i       v       p   '     ������� � ������������'               t � t � 
2    v 8 x ,         >  tm       v      p   '     ������� � ������������'               | � | � 
2    { ; } /       !  �  �p       v      p   '     ������� � ������������'               � � � � 
2    � > � 2       *  j  |t       v      p   '    ������� � ������������'               � � � � 
2    � A � 5       3      x       v      p   '    ������� � ������������'               � � � � 
2    � D � 8       <  �  �{       v      p   '    ������� � ������������'               � � � � 
2    � G � ;       E  ,         v      p   '    ������� � ������������'               � � � � 
2    � J � >       N  �  ��       v      p   '    ������� � ������������'               � � � � 
2    � M � A       W  X  �       v      p   '    ������� � ������������'               � � � � 
2    � P � D       `  �  ��       v 	     p   '    ������� � ������������'               � � � � 
2    � < � 0       �  F  �       w       q   (     ������� � ������������(               � � � � 
2    � ? � 3       �  �  ֵ       w      q   (     ������� � ������������(               � � � � 
2    � B � 6       �  �  º       w      q   (     ������� � ������������(               � � � � 
2    � E � 9       �  b  ��       w      q   (    ������� � ������������(               � � � � 
2    � H � <       �    ��       w      q   (    ������� � ������������(               � � � � 
2    � K � ?         �  ��       w      q   (    ������� � ������������(               � � � � 
2    � N � B         ~  r�       w      q   (    ������� � ������������(               � � 
2    � Q � E         2  ^�       w      q   (    ������� � ������������(               � � 
2    � T � H       )  �  J�       w      q   (    ������� � ������������(               � � 
2    � W � K       6  �  6�       w 	     q   (    ������� � ������������(               � � 
2    � B � 6       �  j"  P      x       r   )     ������� � �����  �  )               � � 
2    � F � :       �  <#  �      x      r   )     ������� � �����  �  )               � � 
2    � J � >       �  $  p       x      r   )     ������� � �����  �  )               � #� #
2    � N � B       �  �$   '      x      r   )    ������� � �����  �  )               ..
2    � R � F         �%  �-      x      r   )    ������� � �����  �  )               99
2    � V � J         �&   4      x      r   )    ������� � �����  �  )               DD
2    � Z � N       %  V'  �:      x      r   )    ������� � �����  �  )               %O%O
2    � ^ � R       6  ((  @A      x      r   )    ������� � �����  �  )               0Z0Z
2    � b � V       G  �(  �G      x      r   )    ������� � �����  �  )               ;e;e
2    � f � Z       X  �)  `N      x 	     r   )    ������� � �����  �  )              ��    2    &             	      �        �       �   *     ���������� ������������*              ��    2    *                >  |        �      �   *     ���������� ������������*              ��    2    .                \  �        �      �   *     ���������� ������������*              ��   	 2    2                z  �        �      �   *    ���������� ������������*              ��  	  2    6                �  0        �      �   *    ���������� ������������*              ��    2    :                �  l        �      �   *    ���������� ������������*              ��    2    >                �  �        �      �   *    ���������� ������������*              ��     2    B                �  �        �      �   *    ���������� ������������*              ��  "   2    F                           �      �   *    ���������� ������������*              ��" $   2    J                .  \        � 	     �   *    ���������� ������������*              �� "   2    7 2           #   �  �        �       �   +     ���������� ������������+              ��# &   2    ; 6           %   �  �        �      �   +     ���������� ������������+              ��' *   2    ? :           '     Z        �      �   +     ���������� ������������+              ��+ .   2    C >           )   Z          �      �   +    ���������� ������������+              ��/ 2   2    G B           *   �  �        �      �   +    ���������� ������������+              ��3 6  " 2    K F           ,   �  v        �      �   +    ���������� ������������+              ��7 : " % 2    O J           .     *        �      �   +    ���������� ������������+              ��; > % ( 2    S N           0   J  �        �      �   +    ���������� ������������+              ��? B ( + 2    W R           2   �  �        �      �   +    ���������� ������������+              ��C F + . 2    [ V           3   �  F        � 	     �   +    ���������� ������������+              ��< @ # ' 2    H C          N   �  �        �       �   ,     ���������� ������������,              ��A F ' , 2    M H !         R     0         �      �   ,     ���������� ������������,              ��F L + 1 2    R M $         V   f  �!        �      �   ,     ���������� ������������,              ��K R / 6 2    W R '         Y   �   #        �      �   ,    ���������� ������������,              ��P X 3 ; 2    \ W *         ]   	  h$        �      �   ,    ���������� ������������,              ��U ^ 7 @ 2    a \ -         `   t	  �%        �      �   ,    ���������� ������������,              ��Z d ; E 2    f a 0         d   �	  8'        �      �   ,    ���������� ������������,              ��_ j ? J 2    k f 3         h   (
  �(        �      �   ,    ���������� ������������,              ��d p C O 2    p k 6         k   �
  *        �      �   ,    ���������� ������������,              ��i v G T 2    u p 9         o   �
  p+        � 	     �   ,    ���������� ������������,              ��] m : J 2    b ] &        �   D  T=        �       �   -     ���������� ������������-              ��d u @ P 2    g b )        �   �  �?        �      �   -     ���������� ������������-              ��k } F V 2    l g ,         �   4  B        �      �   -     ���������� ������������-              ��r � L \ 2    q l / #       �   �  \D        �      �   -    ���������� ������������-              ��y � R b 2    v q 2 &       �   $  �F        �      �   -    ���������� ������������-              ��� � X h 2    { v 5 )       �   �  I        �      �   -    ���������� ������������-              ��� � ^ n 2    � { 8 ,       �     dK        �      �   -    ���������� ������������-              ��� � d t 2    � � ; /       �   �  �M        �      �   -    ���������� ������������-              ��� � j z 2    � � > 2       �     P        �      �   -    ���������� ������������-              ��� � p � 2    � � A 5       �   |  lR        � 	     �   -    ���������� ������������-              ��� � _ q 2    { v - !         \  (n        �       �   .     ���������� ������������.              ��� � f y 2    � { 0 $       #  �  �q        �      �   .     ���������� ������������.              ��� � m � 2    � � 3 '       ,  �  0u        �      �   .     ���������� ������������.              ��� � t � 2    � � 6 *       5    �x        �      �   .    ���������� ������������.              ��� � { � 2    � � 9 -       >  �  8|        �      �   .    ���������� ������������.              ��� � � � 2    � � < 0       G  J  �        �      �   .    ���������� ������������.              ��� � � � 2    � � ? 3       P  �  @�        �      �   .    ���������� ������������.              ��� � � � 2    � � B 6       Y  v  Ć        �      �   .    ���������� ������������.              ��� � � � 2    � � E 9       b    H�        �      �   .    ���������� ������������.              ��� � � � 2    � � H <       k  �  ̍        � 	     �   .    ���������� ������������.              ��� � � � 2    � � 4 (       �  �  ֵ        �       �   /     ���������� ������������/              ��� � � � 2    � � 7 +       �  �  º        �      �   /     ���������� ������������/              ��� � � � 2    � � : .       �  b  ��        �      �   /     ���������� ������������/              ��� 	� � 2    � � = 1       �    ��        �      �   /    ���������� ������������/              ��� � � 2    � � @ 4         �  ��        �      �   /    ���������� ������������/              ��� � � 2    � � C 7         ~  r�        �      �   /    ���������� ������������/              ��*� � 2    � � F :         2  ^�        �      �   /    ���������� ������������/              ��5� � 2    � � I =       )  �  J�        �      �   /    ���������� ������������/              ��@� � 2    � � L @       6  �  6�        �      �   /    ���������� ������������/              ��$K� � 2    � � O C       B  N   "�        � 	     �   /    ���������� ������������/              ��6� � 2    � � : .       �  #  �       �       �   0     ���������� �����  �  0              ��C� � 2    � � > 2       �  �#  �       �      �   0     ���������� �����  �  0              ��$P� � 2    � � B 6       �  �$  &       �      �   0     ���������� �����  �  0              ��0]� � 2    � � F :         �%  �,       �      �   0    ���������� �����  �  0              ��<j� 	2    � � J >         f&  03       �      �   0    ���������� �����  �  0              ��Hw� 2    � � N B       #  8'  �9       �      �   0    ���������� �����  �  0              ��T�� 2    � � R F       4  
(  P@       �      �   0    ���������� �����  �  0              ��`�� '2    � � V J       D  �(  �F       �      �   0    ���������� �����  �  0              ��l�12    � � Z N       U  �)  pM       �      �   0    ���������� �����  �  0              ��x�;2    � � ^ R       f  �*   T       � 	     �   0    ���������� �����  �  0           ����              6             	      �               ��1         ���� � ������������1           ����              ;                >  |              ��1         ���� � ������������1           ����   	 
          @                \  �              ��1         ���� � ������������1           ����              E                z  �              ��1        ���� � ������������1           ����              J                �  0              ��1        ���� � ������������1           ����              O                �  l              ��1        ���� � ������������1           ����              T                �  �              ��1        ���� � ������������1           ����              Y                �  �              ��1        ���� � ������������1           ����              ^                                 ��1        ���� � ������������1           ����              c                .  \       	       ��1        ���� � ������������1           ����   
           Q $           #   �  �               ��2         ���� � ������������2           ����              V (           %   �  �              ��2         ���� � ������������2           ����              [ ,           '     Z              ��2         ���� � ������������2           ����              ` 0           )   Z                ��2        ���� � ������������2           ����              e 4           *   �  �              ��2        ���� � ������������2           ����              j 8           ,   �  v              ��2        ���� � ������������2           ����              o <           .     *              ��2        ���� � ������������2           ����              t @           0   J  �              ��2        ���� � ������������2           ����              y D           2   �  �              ��2        ���� � ������������2           ����              ~ H           3   �  F       	       ��2        ���� � ������������2           ����              k 5          N   �  �               ��3         ���� � ������������3          ����              p 9 !         R     0               ��3         ���� � ������������3          ����              u = $         V   f  �!              ��3         ���� � ������������3          ����              z A '         Y   �   #              ��3        ���� � ������������3          ����               E *         ]   	  h$              ��3        ���� � ������������3          ����              � I -         `   t	  �%              ��3        ���� � ������������3          ����              � M 0         d   �	  8'              ��3        ���� � ������������3          ����              � Q 3         h   (
  �(              ��3        ���� � ������������3          ����   ! "          � U 6         k   �
  *              ��3        ���� � ������������3          ����   # $          � Y 9         o   �
  p+       	       ��3        ���� � ������������3           ����              � E &        �   D  T=               ��4         ���� � ������������4          ����              � I )        �   �  �?              ��4         ���� � ������������4          ����              � M ,         �   4  B              ��4         ���� � ������������4          ����              � Q / #       �   �  \D              ��4        ���� � ������������4          ����              � U 2 &       �   $  �F              ��4        ���� � ������������4          ����               � Y 5 )       �   �  I              ��4        ���� � ������������4          ����   ! "          � ] 8 ,       �     dK              ��4        ���� � ������������4          ����   # $          � a ; /       �   �  �M              ��4        ���� � ������������4          ����   & '          � e > 2       �     P              ��4        ���� � ������������4          ����   ( )          � i A 5       �   |  lR       	       ��4        ���� � ������������4           ����              + . /         	      �       *        ��5         ���� � ������������5           ����              - 1 4            >  |       *       ��5         ���� � ������������5           ����              / 4 9            \  �       *       ��5         ���� � ������������5           ����   	 
          1 7 >            z  �       *       ��5        ���� � ������������5           ����              3 : C            �  0       *       ��5        ���� � ������������5           ����              5 = H            �  l       *       ��5        ���� � ������������5           ����              7 @ M            �  �       *       ��5        ���� � ������������5           ����              9 C R            �  �       *       ��5        ���� � ������������5           ����              ; F W                      *       ��5        ���� � ������������5           ����              = I \            .  \       *	       ��5        ���� � ������������5           ����              * 6 J        #   �  �       +        ��6         ���� � ������������6           ����   	 
          - 9 O        %   �  �       +       ��6         ���� � ������������6           ����              0 < T        '     Z       +       ��6         ���� � ������������6           ����              3 ? Y        )   Z         +       ��6        ���� � ������������6           ����              6 B ^        *   �  �       +       ��6        ���� � ������������6           ����              9 E c        ,   �  v       +       ��6        ���� � ������������6           ����              < H h         .     *       +       ��6        ���� � ������������6           ����              ? K m "       0   J  �       +       ��6        ���� � ������������6           ����              B N r $       2   �  �       +       ��6        ���� � ������������6           ����              E Q w &       3   �  F       +	       ��6        ���� � ������������6           ����              2 = d        N   �  �       ,        ��7         ���� � ������������7          ����              5 A i        R     0        ,       ��7         ���� � ������������7          ����              8 E n        V   f  �!       ,       ��7         ���� � ������������7          ����              ; I s !       Y   �   #       ,       ��7        ���� � ������������7          ����              > M x $       ]   	  h$       ,       ��7        ���� � ������������7          ����              A Q } '       `   t	  �%       ,       ��7        ���� � ������������7          ����              D U � *       d   �	  8'       ,       ��7        ���� � ������������7          ����              G Y � -       h   (
  �(       ,       ��7        ���� � ������������7          ����              J ] � 0       k   �
  *       ,       ��7        ���� � ������������7          ����              M a � 3       o   �
  p+       ,	       ��7        ���� � ������������7           ����              : N }         �   D  T=       -        ��8         ���� � ������������8          ����              = R � #       �   �  �?       -       ��8         ���� � ������������8          ����              @ V � &       �   4  B       -       ��8         ���� � ������������8          ����              C Z � )       �   �  \D       -       ��8        ���� � ������������8          ����              F ^ � ,       �   $  �F       -       ��8        ���� � ������������8          ����              I b � /       �   �  I       -       ��8        ���� � ������������8          ����              L f � 2       �     dK       -       ��8        ���� � ������������8          ����              O j � 5       �   �  �M       -       ��8        ���� � ������������8          ����     !          R n � 8       �     P       -       ��8        ���� � ������������8          ����   " #          U r � ;       �   |  lR       -	       ��8        ���� � ������������8           ����             !                ,  h       �        ��9         ���� � ������������9           ����             &                J  �       �       ��9         ���� � ������������9           ����             +                h  �       �       ��9         ���� � ������������9           ����  
           0                �         �       ��9        ���� � ������������9           ����             5                �  H       �       ��9        ���� � ������������9           ����             :             	   �  �       �       ��9        ���� � ������������9           ����             ?             	   �  �       �       ��9        ���� � ������������9           ����             D             
   �  �       �       ��9        ���� � ������������9           ����             I             
     8       �       ��9        ���� � ������������9           ����             N                :  t       �	       ��9        ���� � ������������9           ����   	          < $              �         �        ��:         ���� � ������������:           ����  
           A (              �  �       �       ��:         ���� � ������������:           ����             F ,              *  ~	       �       ��:         ���� � ������������:           ����             K 0              f  2
       �       ��:        ���� � ������������:           ����             P 4              �  �
       �       ��:        ���� � ������������:           ����             U 8              �  �       �       ��:        ���� � ������������:           ����             Z <                N       �       ��:        ���� � ������������:           ����             _ @           !   V         �       ��:        ���� � ������������:           ����             d D           #   �  �       �       ��:        ���� � ������������:           ����             i H           $   �  j       �	       ��:        ���� � ������������:           ����             V 5          :   �  �       �        ��;         ���� � ������������;          ����             [ 9 !         >     `       �       ��;         ���� � ������������;          ����             ` = $         B   r  �       �       ��;         ���� � ������������;          ����             e A '         E   �  0       �       ��;        ���� � ������������;          ����             j E *         I   &  �       �       ��;        ���� � ������������;          ����             o I -         L   �          �       ��;        ���� � ������������;          ����             t M 0         P   �  h       �       ��;        ���� � ������������;          ����             y Q 3         T   4  �        �       ��;        ���� � ������������;          ����              ~ U 6         W   �  8"       �       ��;        ���� � ������������;          ����  ! "          � Y 9         [   �  �#       �	       ��;        ���� � ������������;           ����             o E &        �   P
  �3       �        ��<         ���� � ������������<          ����             u I )        �   �
  �5       �       ��<         ���� � ������������<          ����             { M ,         �   @  @8       �       ��<         ���� � ������������<          ����             � Q / #       �   �  �:       �       ��<        ���� � ������������<          ����             � U 2 &       �   0  �<       �       ��<        ���� � ������������<          ����             � Y 5 )       �   �  H?       �       ��<        ���� � ������������<          ����              � ] 8 ,       �      �A       �       ��<        ���� � ������������<          ����  ! "          � a ; /       �   �  �C       �       ��<        ���� � ������������<          ����  $ %          � e > 2       �     PF       �       ��<        ���� � ������������<          ����  & '          � i A 5       �   �  �H       �	       ��<        ���� � ������������<           ����                           ,  h       �        ��=         ���� � ������������=           ����                           J  �       �       ��=         ���� � ������������=           ����               $            h  �       �       ��=         ���� � ������������=           ����   	           " )            �         �       ��=        ���� � ������������=           ����  
            % .            �  H       �       ��=        ���� � ������������=           ����               ( 3         	   �  �       �       ��=        ���� � ������������=           ����             " + 8         	   �  �       �       ��=        ���� � ������������=           ����             $ . =         
   �  �       �       ��=        ���� � ������������=           ����             & 1 B         
     8       �       ��=        ���� � ������������=           ����             ( 4 G            :  t       �	       ��=        ���� � ������������=           ����              ! 5           �         �        ��>         ���� � ������������>           ����   	           $ :           �  �       �       ��>         ���� � ������������>           ����  
            ' ?           *  ~	       �       ��>         ���� � ������������>           ����              * D           f  2
       �       ��>        ���� � ������������>           ����             ! - I           �  �
       �       ��>        ���� � ������������>           ����             $ 0 N           �  �       �       ��>        ���� � ������������>           ����             ' 3 S              N       �       ��>        ���� � ������������>           ����             * 6 X "       !   V         �       ��>        ���� � ������������>           ����             - 9 ] $       #   �  �       �       ��>        ���� � ������������>           ����             0 < b &       $   �  j       �	       ��>        ���� � ������������>           ����  
            ( O        :   �  �       �        ��?         ���� � ������������?          ����               , T        >     `       �       ��?         ���� � ������������?          ����             # 0 Y        B   r  �       �       ��?         ���� � ������������?          ����             & 4 ^ !       E   �  0       �       ��?        ���� � ������������?          ����             ) 8 c $       I   &  �       �       ��?        ���� � ������������?          ����             , < h '       L   �          �       ��?        ���� � ������������?          ����             / @ m *       P   �  h       �       ��?        ���� � ������������?          ����             2 D r -       T   4  �        �       ��?        ���� � ������������?          ����             5 H w 0       W   �  8"       �       ��?        ���� � ������������?          ����             8 L | 3       [   �  �#       �	       ��?        ���� � ������������?           ����             % 9 h         �   P
  �3       �        ��@         ���� � ������������@          ����             ( = n #       �   �
  �5       �       ��@         ���� � ������������@          ����             + A t &       �   @  @8       �       ��@         ���� � ������������@          ����             . E z )       �   �  �:       �       ��@        ���� � ������������@          ����             1 I � ,       �   0  �<       �       ��@        ���� � ������������@          ����             4 M � /       �   �  H?       �       ��@        ���� � ������������@          ����             7 Q � 2       �      �A       �       ��@        ���� � ������������@          ����             : U � 5       �   �  �C       �       ��@        ���� � ������������@          ����              = Y � 8       �     PF       �       ��@        ���� � ������������@          ����  ! "          @ ] � ;       �   �  �H       �	       ��@        ���� � ������������@             ��              H            �����
  �         �       �    A         ���� � ������������A             ��   	           M            ����          �      �    A         ���� � ������������A             ��  
            R            ����,  X        �      �    A         ���� � ������������A             ��              W            ����J  �        �      �    A         ���� � ������������A             ��              \            ����h  �        �      �    A         ���� � ������������A             ��              a            �����          �      �    A         ���� � ������������A             ��              f            �����  H        �      �    A         ���� � ������������A             ��              k            �����  �        �      �    A         ���� � ������������A             ��              p            �����  �        �      �    A         ���� � ������������A             ��              u            �����  �        � 	     �    A         ���� � ������������A            ��              c $     (     ����v  b%        �       �    B         ���� � ������������B            ��              h (     (     �����  &        �      �    B         ���� � ������������B            ��              m ,     (     �����  �&        �      �    B         ���� � ������������B            ��              r 0     (     ����*  ~'        �      �    B         ���� � ������������B            ��              w 4     (     ����f  2(        �      �    B         ���� � ������������B            ��              | 8     (     �����  �(        �      �    B         ���� � ������������B            ��              � <     (     �����  �)        �      �    B         ���� � ������������B            ��              � @     (     ����  N*        �      �    B         ���� � ������������B            ��              � D     (     ����V  +        �      �    B         ���� � ������������B            ��               � H     (     �����  �+        � 	     �    B         ���� � ������������B           ��              } 5    2     �����  >        �       �    C         ���� � ������������C           ��              � 9 !   2     �����  p?        �      �    C         ���� � ������������C           ��              � = $   2     ����6  �@        �      �    C         ���� � ������������C           ��              � A '   2     �����  @B        �      �    C         ���� � ������������C           ��              � E *   2     �����  �C        �      �    C         ���� � ������������C           ��              � I -   2     ����D  E        �      �    C         ���� � ������������C           ��              � M 0   2     �����  xF        �      �    C         ���� � ������������C           ��               � Q 3   2     �����  �G        �      �    C         ���� � ������������C           ��  " #           � U 6   2     ����R  HI        �      �    C         ���� � ������������C           ��  $ %           � Y 9   2     �����  �J        � 	     �    C         ���� � ������������C          	 ��              � E &  <     ����  dd        �       �    D         ���� � ������������D          	 ��              � I )  <     �����  �f        �      �    D         ���� � ������������D          	 ��              � M ,   <     ����  i        �      �    D         ���� � ������������D          	 ��              � Q / # <     ����|  lk        �      �    D         ���� � ������������D          	 ��              � U 2 & <     �����  �m        �      �    D         ���� � ������������D          	 ��    !           � Y 5 ) <     ����l  p        �      �    D         ���� � ������������D          	 ��  " #           � ] 8 , <     �����  tr        �      �    D         ���� � ������������D          	 ��  $ %           � a ; / <     ����\  �t        �      �    D         ���� � ������������D          	 ��  ' (           � e > 2 <     �����  $w        �      �    D         ���� � ������������D          	 ��  ) *           � i A 5 <     ����L  |y        � 	     �    D         ���� � ������������D             ��              < @ A        �����
  �         �       �    E         ���� � ������������E             ��              > C F        ����          �      �    E         ���� � ������������E             ��              @ F K        ����,  X        �      �    E         ���� � ������������E             ��  	 
           B I P        ����J  �        �      �    E         ���� � ������������E             ��              D L U        ����h  �        �      �    E         ���� � ������������E             ��              F O Z        �����          �      �    E         ���� � ������������E             ��              H R _        �����  H        �      �    E         ���� � ������������E             ��              J U d        �����  �        �      �    E         ���� � ������������E             ��              L X i        �����  �        �      �    E         ���� � ������������E             ��              N [ n        �����  �        � 	     �    E         ���� � ������������E            ��              ; H \  (     ����v  b%        �       �    F         ���� � ������������F            ��  	 
           > K a  (     �����  &        �      �    F         ���� � ������������F            ��              A N f  (     �����  �&        �      �    F         ���� � ������������F            ��              D Q k  (     ����*  ~'        �      �    F         ���� � ������������F            ��              G T p  (     ����f  2(        �      �    F         ���� � ������������F            ��              J W u  (     �����  �(        �      �    F         ���� � ������������F            ��              M Z z   (     �����  �)        �      �    F         ���� � ������������F            ��              P ]  " (     ����  N*        �      �    F         ���� � ������������F            ��              S ` � $ (     ����V  +        �      �    F         ���� � ������������F            ��              V c � & (     �����  �+        � 	     �    F         ���� � ������������F           ��              C O v  2     �����  >        �       �    G         ���� � ������������G           ��              F S {  2     �����  p?        �      �    G         ���� � ������������G           ��              I W �  2     ����6  �@        �      �    G         ���� � ������������G           ��              L [ � ! 2     �����  @B        �      �    G         ���� � ������������G           ��              O _ � $ 2     �����  �C        �      �    G         ���� � ������������G           ��              R c � ' 2     ����D  E        �      �    G         ���� � ������������G           ��              U g � * 2     �����  xF        �      �    G         ���� � ������������G           ��              X k � - 2     �����  �G        �      �    G         ���� � ������������G           ��              [ o � 0 2     ����R  HI        �      �    G         ���� � ������������G           ��              ^ s � 3 2     �����  �J        � 	     �    G         ���� � ������������G          	 ��              K ` �   <     ����  dd        �       �    H         ���� � ������������H          	 ��              N d � # <     �����  �f        �      �    H         ���� � ������������H          	 ��              Q h � & <     ����  i        �      �    H         ���� � ������������H          	 ��              T l � ) <     ����|  lk        �      �    H         ���� � ������������H          	 ��              W p � , <     �����  �m        �      �    H         ���� � ������������H          	 ��              Z t � / <     ����l  p        �      �    H         ���� � ������������H          	 ��              ] x � 2 <     �����  tr        �      �    H         ���� � ������������H          	 ��              ` | � 5 <     ����\  �t        �      �    H         ���� � ������������H          	 ��    !           c � � 8 <     �����  $w        �      �    H         ���� � ������������H          	 ��  " #           f � � ; <     ����L  |y        � 	     �    H         ���� � ������������H           ����             .                �   �        �        ��I         ���� � ������������I           ����             3                �   �       �       ��I         ���� � ������������I           ����   	          8                         �       ��I         ���� � ������������I           ����             =                "  D       �       ��I        ���� � ������������I           ����             B                @  �       �       ��I        ���� � ������������I           ����             G                ^  �       �       ��I        ���� � ������������I           ����             L                |  �       �       ��I        ���� � ������������I           ����             Q                �  4       �       ��I        ���� � ������������I           ����             V                �  p       �       ��I        ���� � ������������I           ����             [             	   �  �       �	       ��I        ���� � ������������I           ����  	 
          I $              N  �       �        ��J         ���� � ������������J           ����             N (              �  �       �       ��J         ���� � ������������J           ����             S ,              �  R       �       ��J         ���� � ������������J           ����             X 0                	       �       ��J        ���� � ������������J           ����             ] 4              >  �	       �       ��J        ���� � ������������J           ����             b 8              z  n
       �       ��J        ���� � ������������J           ����             g <              �  "       �       ��J        ���� � ������������J           ����             l @              �  �       �       ��J        ���� � ������������J           ����             q D               .  �       �       ��J        ���� � ������������J           ����             v H           !   j  >       �	       ��J        ���� � ������������J          ����             c 5          6   Z  h       �        ��K         ���� � ������������K          ����             h 9 !         :   �  �       �       ��K         ���� � ������������K          ����             m = $         >     8       �       ��K         ���� � ������������K          ����             r A '         A   h  �       �       ��K        ���� � ������������K          ����             w E *         E   �         �       ��K        ���� � ������������K          ����             | I -         H     p       �       ��K        ���� � ������������K          ����             � M 0         L   v  �       �       ��K        ���� � ������������K          ����             � Q 3         P   �  @       �       ��K        ���� � ������������K          ����    !          � U 6         S   *  �        �       ��K        ���� � ������������K          ����  " #          � Y 9         W   �  "       �	       ��K        ���� � ������������K          ����             | E &           �	  �1       �        ��L         ���� � ������������L          ����             � I )        �   d
  �3       �       ��L         ���� � ������������L          ����             � M ,         �   �
  L6       �       ��L         ���� � ������������L          ����             � Q / #       �   T  �8       �       ��L        ���� � ������������L          ����             � U 2 &       �   �  �:       �       ��L        ���� � ������������L          ����             � Y 5 )       �   D  T=       �       ��L        ���� � ������������L          ����    !          � ] 8 ,       �   �  �?       �       ��L        ���� � ������������L          ����  " #          � a ; /       �   4  B       �       ��L        ���� � ������������L          ����  % &          � e > 2       �   �  \D       �       ��L        ���� � ������������L          ����  ' (          � i A 5       �   $  �F       �	       ��L        ���� � ������������L           ����             # & '            �   �                ��M         ���� � ������������M           ����             % ) ,            �   �              ��M         ���� � ������������M           ����             ' , 1                            ��M         ���� � ������������M           ����   	          ) / 6            "  D              ��M        ���� � ������������M           ����  
           + 2 ;            @  �              ��M        ���� � ������������M           ����             - 5 @            ^  �              ��M        ���� � ������������M           ����             / 8 E            |  �              ��M        ���� � ������������M           ����             1 ; J            �  4              ��M        ���� � ������������M           ����             3 > O            �  p              ��M        ���� � ������������M           ����             5 A T         	   �  �       	       ��M        ���� � ������������M           ����             " . B           N  �               ��N         ���� � ������������N           ����   	          % 1 G           �  �              ��N         ���� � ������������N           ����  
           ( 4 L           �  R              ��N         ���� � ������������N           ����             + 7 Q             	              ��N        ���� � ������������N           ����             . : V           >  �	              ��N        ���� � ������������N           ����             1 = [           z  n
              ��N        ���� � ������������N           ����             4 @ `            �  "              ��N        ���� � ������������N           ����             7 C e "          �  �              ��N        ���� � ������������N           ����             : F j $           .  �              ��N        ���� � ������������N           ����             = I o &       !   j  >       	       ��N        ���� � ������������N          ����  
           * 5 \        6   Z  h               ��O         ���� � ������������O          ����             - 9 a        :   �  �              ��O         ���� � ������������O          ����             0 = f        >     8              ��O         ���� � ������������O          ����             3 A k !       A   h  �              ��O        ���� � ������������O          ����             6 E p $       E   �                ��O        ���� � ������������O          ����             9 I u '       H     p              ��O        ���� � ������������O          ����             < M z *       L   v  �              ��O        ���� � ������������O          ����             ? Q  -       P   �  @              ��O        ���� � ������������O          ����             B U � 0       S   *  �               ��O        ���� � ������������O          ����             E Y � 3       W   �  "       	       ��O        ���� � ������������O          ����             2 F u            �	  �1               ��P         ���� � ������������P          ����             5 J { #       �   d
  �3              ��P         ���� � ������������P          ����             8 N � &       �   �
  L6              ��P         ���� � ������������P          ����             ; R � )       �   T  �8              ��P        ���� � ������������P          ����             > V � ,       �   �  �:              ��P        ���� � ������������P          ����             A Z � /       �   D  T=              ��P        ���� � ������������P          ����             D ^ � 2       �   �  �?              ��P        ���� � ������������P          ����             G b � 5       �   4  B              ��P        ���� � ������������P          ����              J f � 8       �   �  \D              ��P        ���� � ������������P          ����  ! "          M j � ;       �   $  �F       	       ��P        ���� � ������������P           ����                          !   �  /       V        ��Q         ���� � ������������Q           ����             !             (   �  �       V       ��Q         ���� � ������������Q           ����             &             )            V       ��Q         ���� � ������������Q           ����  
           +             )   *  T       V       ��Q        ���� � ������������Q           ����             0             *   H  �       V       ��Q        ���� � ������������Q           ����             5             +   f  �       V       ��Q        ���� � ������������Q           ����             :             +   �         V       ��Q        ���� � ������������Q           ����             ?             ,   �  D       V       ��Q        ���� � ������������Q           ����             D             ,   �  �       V       ��Q        ���� � ������������Q           ����             I             -   �  �       V	       ��Q        ���� � ������������Q           ����   	          7 $           G   V	         W        ��R         ���� � ������������R           ����  
           < (           I   �	  �       W       ��R         ���� � ������������R           ����             A ,           K   �	  j       W       ��R         ���� � ������������R           ����             F 0           M   

         W       ��R        ���� � ������������R           ����             K 4           N   F
  �       W       ��R        ���� � ������������R           ����             P 8           P   �
  �       W       ��R        ���� � ������������R           ����             U <           R   �
  :        W       ��R        ���� � ������������R           ����             Z @           T   �
  �        W       ��R        ���� � ������������R           ����             _ D           V   6  �!       W       ��R        ���� � ������������R           ����             d H           W   r  V"       W	       ��R        ���� � ������������R           ����             Q 5          ~   b  �1       X        ��S         ���� � ������������S          ����             V 9 !         �   �  �2       X       ��S         ���� � ������������S          ����             [ = $         �     X4       X       ��S         ���� � ������������S          ����             ` A '         �   p  �5       X       ��S        ���� � ������������S          ����             e E *         �   �  (7       X       ��S        ���� � ������������S          ����             j I -         �   $  �8       X       ��S        ���� � ������������S          ����             o M 0         �   ~  �9       X       ��S        ���� � ������������S          ����             t Q 3         �   �  `;       X       ��S        ���� � ������������S          ����              y U 6         �   2  �<       X       ��S        ���� � ������������S          ����  ! "          ~ Y 9         �   �  0>       X	       ��S        ���� � ������������S           ����             j E &        �   �  �T       Y        ��T         ���� � ������������T          ����             p I )        �   l  W       Y       ��T         ���� � ������������T          ����             v M ,         �   �  tY       Y       ��T         ���� � ������������T          ����             | Q / #       �   \  �[       Y       ��T        ���� � ������������T          ����             � U 2 &       �   �  $^       Y       ��T        ���� � ������������T          ����             � Y 5 )       �   L  |`       Y       ��T        ���� � ������������T          ����              � ] 8 ,       �   �  �b       Y       ��T        ���� � ������������T          ����  ! "          � a ; /         <  ,e       Y       ��T        ���� � ������������T          ����  $ %          � e > 2       	  �  �g       Y       ��T        ���� � ������������T          ����  & '          � i A 5         ,  �i       Y	       ��T        ���� � ������������T           ����                        !   �  /       g        ��U         ���� � ������������U           ����                        (   �  �       g       ��U         ���� � ������������U           ����                        )            g       ��U         ���� � ������������U           ����   	            $         )   *  T       g       ��U        ���� � ������������U           ����  
              )         *   H  �       g       ��U        ���� � ������������U           ����              # .         +   f  �       g       ��U        ���� � ������������U           ����              & 3         +   �         g       ��U        ���� � ������������U           ����              ) 8         ,   �  D       g       ��U        ���� � ������������U           ����             ! , =         ,   �  �       g       ��U        ���� � ������������U           ����             # / B         -   �  �       g	       ��U        ���� � ������������U           ����               0        G   V	         h        ��V         ���� � ������������V           ����   	            5        I   �	  �       h       ��V         ���� � ������������V           ����  
            " :        K   �	  j       h       ��V         ���� � ������������V           ����              % ?        M   

         h       ��V        ���� � ������������V           ����              ( D        N   F
  �       h       ��V        ���� � ������������V           ����              + I        P   �
  �       h       ��V        ���� � ������������V           ����             " . N         R   �
  :        h       ��V        ���� � ������������V           ����             % 1 S "       T   �
  �        h       ��V        ���� � ������������V           ����             ( 4 X $       V   6  �!       h       ��V        ���� � ������������V           ����             + 7 ] &       W   r  V"       h	       ��V        ���� � ������������V           ����  
            # J        ~   b  �1       i        ��W         ���� � ������������W          ����              ' O        �   �  �2       i       ��W         ���� � ������������W          ����              + T        �     X4       i       ��W         ���� � ������������W          ����             ! / Y !       �   p  �5       i       ��W        ���� � ������������W          ����             $ 3 ^ $       �   �  (7       i       ��W        ���� � ������������W          ����             ' 7 c '       �   $  �8       i       ��W        ���� � ������������W          ����             * ; h *       �   ~  �9       i       ��W        ���� � ������������W          ����             - ? m -       �   �  `;       i       ��W        ���� � ������������W          ����             0 C r 0       �   2  �<       i       ��W        ���� � ������������W          ����             3 G w 3       �   �  0>       i	       ��W        ���� � ������������W           ����               4 c         �   �  �T       j        ��X         ���� � ������������X          ����             # 8 i #       �   l  W       j       ��X         ���� � ������������X          ����             & < o &       �   �  tY       j       ��X         ���� � ������������X          ����             ) @ u )       �   \  �[       j       ��X        ���� � ������������X          ����             , D { ,       �   �  $^       j       ��X        ���� � ������������X          ����             / H � /       �   L  |`       j       ��X        ���� � ������������X          ����             2 L � 2       �   �  �b       j       ��X        ���� � ������������X          ����             5 P � 5         <  ,e       j       ��X        ���� � ������������X          ����              8 T � 8       	  �  �g       j       ��X        ���� � ������������X          ����  ! "          ; X � ;         ,  �i       j	       ��X        ���� � ������������X           ����             C                @  �       �         ��Y         ���� � ������������Y           ����   	          H                 ^  �       �        ��Y         ���� � ������������Y           ����  
           M             !   |  �       �        ��Y         ���� � ������������Y           ����             R             !   �  4       �        ��Y        ���� � ������������Y           ����             W             "   �  p       �        ��Y        ���� � ������������Y           ����             \             #   �  �       �        ��Y        ���� � ������������Y           ����             a             #   �  �       �        ��Y        ���� � ������������Y           ����             f             $     $       �        ��Y        ���� � ������������Y           ����             k             $   0  `       �        ��Y        ���� � ������������Y           ����             p             %   N  �       �	        ��Y        ���� � ������������Y           ����             ^ $           ;   �  R       �        ��Z         ���� � ������������Z           ����             c (           =            �       ��Z         ���� � ������������Z           ����             h ,           ?   >  �       �       ��Z         ���� � ������������Z           ����             m 0           A   z  n       �       ��Z        ���� � ������������Z           ����             r 4           B   �  "       �       ��Z        ���� � ������������Z           ����             w 8           D   �  �       �       ��Z        ���� � ������������Z           ����             | <           F   .	  �       �       ��Z        ���� � ������������Z           ����             � @           H   j	  >       �       ��Z        ���� � ������������Z           ����             � D           J   �	  �       �       ��Z        ���� � ������������Z           ����              � H           K   �	  �       �	       ��Z        ���� � ������������Z          ����             x 5          n   �
  H+       �        ��[         ���� � ������������[          ����             } 9 !         r   ,  �,       �       ��[         ���� � ������������[          ����             � = $         v   �  .       �       ��[         ���� � ������������[          ����             � A '         y   �  �/       �       ��[        ���� � ������������[          ����             � E *         }   :  �0       �       ��[        ���� � ������������[          ����             � I -         �   �  P2       �       ��[        ���� � ������������[          ����             � M 0         �   �  �3       �       ��[        ���� � ������������[          ����              � Q 3         �   H   5       �       ��[        ���� � ������������[          ����  " #          � U 6         �   �  �6       �       ��[        ���� � ������������[          ����  $ %          � Y 9         �   �  �7       �	       ��[        ���� � ������������[          ����             � E &        �   d  �L       �        ��\         ���� � ������������\          ����             � I )        �   �  LO       �       ��\         ���� � ������������\          ����             � M ,         �   T  �Q       �       ��\         ���� � ������������\          ����             � Q / #       �   �  �S       �       ��\        ���� � ������������\          ����             � U 2 &       �   D  TV       �       ��\        ���� � ������������\          ����    !          � Y 5 )       �   �  �X       �       ��\        ���� � ������������\          ����  " #          � ] 8 ,       �   4  [       �       ��\        ���� � ������������\          ����  $ %          � a ; /       �   �  \]       �       ��\        ���� � ������������\          ����  ' (          � e > 2       �   $  �_       �       ��\        ���� � ������������\          ����  ) *          � i A 5       �   �  b       �	       ��\        ���� � ������������\           ����             7 ; <            @  �       �         ��]         ���� � ������������]           ����             9 > A             ^  �       �        ��]         ���� � ������������]           ����             ; A F         !   |  �       �        ��]         ���� � ������������]           ����  	 
          = D K         !   �  4       �        ��]        ���� � ������������]           ����             ? G P         "   �  p       �        ��]        ���� � ������������]           ����             A J U         #   �  �       �        ��]        ���� � ������������]           ����             C M Z         #   �  �       �        ��]        ���� � ������������]           ����             E P _         $     $       �        ��]        ���� � ������������]           ����             G S d         $   0  `       �        ��]        ���� � ������������]           ����             I V i         %   N  �       �	        ��]        ���� � ������������]           ����             6 C W        ;   �  R       �        ��^         ���� � ������������^           ����  	 
          9 F \        =            �       ��^         ���� � ������������^           ����             < I a        ?   >  �       �       ��^         ���� � ������������^           ����             ? L f        A   z  n       �       ��^        ���� � ������������^           ����             B O k        B   �  "       �       ��^        ���� � ������������^           ����             E R p        D   �  �       �       ��^        ���� � ������������^           ����             H U u         F   .	  �       �       ��^        ���� � ������������^           ����             K X z "       H   j	  >       �       ��^        ���� � ������������^           ����             N [  $       J   �	  �       �       ��^        ���� � ������������^           ����             Q ^ � &       K   �	  �       �	       ��^        ���� � ������������^          ����             > J q        n   �
  H+       �        ��_         ���� � ������������_          ����             A N v        r   ,  �,       �       ��_         ���� � ������������_          ����             D R {        v   �  .       �       ��_         ���� � ������������_          ����             G V � !       y   �  �/       �       ��_        ���� � ������������_          ����             J Z � $       }   :  �0       �       ��_        ���� � ������������_          ����             M ^ � '       �   �  P2       �       ��_        ���� � ������������_          ����             P b � *       �   �  �3       �       ��_        ���� � ������������_          ����             S f � -       �   H   5       �       ��_        ���� � ������������_          ����             V j � 0       �   �  �6       �       ��_        ���� � ������������_          ����             Y n � 3       �   �  �7       �	       ��_        ���� � ������������_          ����             F [ �         �   d  �L       �        ��`         ���� � ������������`          ����             I _ � #       �   �  LO       �       ��`         ���� � ������������`          ����             L c � &       �   T  �Q       �       ��`         ���� � ������������`          ����             O g � )       �   �  �S       �       ��`        ���� � ������������`          ����             R k � ,       �   D  TV       �       ��`        ���� � ������������`          ����             U o � /       �   �  �X       �       ��`        ���� � ������������`          ����             X s � 2       �   4  [       �       ��`        ���� � ������������`          ����             [ w � 5       �   �  \]       �       ��`        ���� � ������������`          ����    !          ^ { � 8       �   $  �_       �       ��`        ���� � ������������`          ����  " #          a  � ;       �   �  b       �	       ��`        ���� � ������������`           ����             )                �  F       "        ��a         ���� � ������������a           ����             .                �  �	       "       ��a         ���� � ������������a           ����   	          3                �  �	       "       ��a         ���� � ������������a           ����             8                
  
       "       ��a        ���� � ������������a           ����             =                (  P
       "       ��a        ���� � ������������a           ����             B                F  �
       "       ��a        ���� � ������������a           ����             G                d  �
       "       ��a        ���� � ������������a           ����             L                �         "       ��a        ���� � ������������a           ����             Q                �  @       "       ��a        ���� � ������������a           ����             V                �  |       "	       ��a        ���� � ������������a           ����  	 
          D $           /   6  �       #        ��b         ���� � ������������b           ����             I (           1   r  V       #       ��b         ���� � ������������b           ����             N ,           3   �  
       #       ��b         ���� � ������������b           ����             S 0           5   �  �       #       ��b        ���� � ������������b           ����             X 4           6   &  r       #       ��b        ���� � ������������b           ����             ] 8           8   b  &       #       ��b        ���� � ������������b           ����             b <           :   �  �       #       ��b        ���� � ������������b           ����             g @           <   �  �       #       ��b        ���� � ������������b           ����             l D           >     B       #       ��b        ���� � ������������b           ����             q H           ?   R  �       #	       ��b        ���� � ������������b           ����             ^ 5          ^   B	  %       $        ��c         ���� � ������������c          ����             c 9 !         b   �	  p&       $       ��c         ���� � ������������c          ����             h = $         f   �	  �'       $       ��c         ���� � ������������c          ����             m A '         i   P
  @)       $       ��c        ���� � ������������c          ����             r E *         m   �
  �*       $       ��c        ���� � ������������c          ����             w I -         p     ,       $       ��c        ���� � ������������c          ����             | M 0         t   ^  x-       $       ��c        ���� � ������������c          ����             � Q 3         x   �  �.       $       ��c        ���� � ������������c          ����    !          � U 6         {     H0       $       ��c        ���� � ������������c          ����  " #          � Y 9            l  �1       $	       ��c        ���� � ������������c           ����             w E &        �   �  $E       %        ��d         ���� � ������������d          ����             } I )        �   L  |G       %       ��d         ���� � ������������d          ����             � M ,         �   �  �I       %       ��d         ���� � ������������d          ����             � Q / #       �   <  ,L       %       ��d        ���� � ������������d          ����             � U 2 &       �   �  �N       %       ��d        ���� � ������������d          ����             � Y 5 )       �   ,  �P       %       ��d        ���� � ������������d          ����    !          � ] 8 ,       �   �  4S       %       ��d        ���� � ������������d          ����  " #          � a ; /       �     �U       %       ��d        ���� � ������������d          ����  % &          � e > 2       �   �  �W       %       ��d        ���� � ������������d          ����  ' (          � i A 5       �     <Z       %	       ��d        ���� � ������������d           ����              ! "            �  F       3        ��e         ���� � ������������e           ����               $ '            �  �	       3       ��e         ���� � ������������e           ����             " ' ,            �  �	       3       ��e         ���� � ������������e           ����   	          $ * 1            
  
       3       ��e        ���� � ������������e           ����  
           & - 6            (  P
       3       ��e        ���� � ������������e           ����             ( 0 ;            F  �
       3       ��e        ���� � ������������e           ����             * 3 @            d  �
       3       ��e        ���� � ������������e           ����             , 6 E            �         3       ��e        ���� � ������������e           ����             . 9 J            �  @       3       ��e        ���� � ������������e           ����             0 < O            �  |       3	       ��e        ���� � ������������e           ����              ) =        /   6  �       4        ��f         ���� � ������������f           ����   	            , B        1   r  V       4       ��f         ���� � ������������f           ����  
           # / G        3   �  
       4       ��f         ���� � ������������f           ����             & 2 L        5   �  �       4       ��f        ���� � ������������f           ����             ) 5 Q        6   &  r       4       ��f        ���� � ������������f           ����             , 8 V        8   b  &       4       ��f        ���� � ������������f           ����             / ; [         :   �  �       4       ��f        ���� � ������������f           ����             2 > ` "       <   �  �       4       ��f        ���� � ������������f           ����             5 A e $       >     B       4       ��f        ���� � ������������f           ����             8 D j &       ?   R  �       4	       ��f        ���� � ������������f           ����  
           % 0 W        ^   B	  %       5        ��g         ���� � ������������g          ����             ( 4 \        b   �	  p&       5       ��g         ���� � ������������g          ����             + 8 a        f   �	  �'       5       ��g         ���� � ������������g          ����             . < f !       i   P
  @)       5       ��g        ���� � ������������g          ����             1 @ k $       m   �
  �*       5       ��g        ���� � ������������g          ����             4 D p '       p     ,       5       ��g        ���� � ������������g          ����             7 H u *       t   ^  x-       5       ��g        ���� � ������������g          ����             : L z -       x   �  �.       5       ��g        ���� � ������������g          ����             = P  0       {     H0       5       ��g        ���� � ������������g          ����             @ T � 3          l  �1       5	       ��g        ���� � ������������g           ����             - A p         �   �  $E       6        ��h         ���� � ������������h          ����             0 E v #       �   L  |G       6       ��h         ���� � ������������h          ����             3 I | &       �   �  �I       6       ��h         ���� � ������������h          ����             6 M � )       �   <  ,L       6       ��h        ���� � ������������h          ����             9 Q � ,       �   �  �N       6       ��h        ���� � ������������h          ����             < U � /       �   ,  �P       6       ��h        ���� � ������������h          ����             ? Y � 2       �   �  4S       6       ��h        ���� � ������������h          ����             B ] � 5       �     �U       6       ��h        ���� � ������������h          ����              E a � 8       �   �  �W       6       ��h        ���� � ������������h          ����  ! "          H e � ;       �     <Z       6	       ��h        ���� � ������������h           ����             ;             2   `	  �       �      �   i         ���� � ������������i           ����             @             0   ~	  �       �     �   i         ���� � ������������i           ����  	 
          E             1   �	  8       �     �   i         ���� � ������������i           ����             J             1   �	  t       �     �   i        ���� � ������������i           ����             O             2   �	  �       �     �   i        ���� � ������������i           ����             T             3   �	  �       �     �   i        ���� � ������������i           ����             Y             3   
  (       �     �   i        ���� � ������������i           ����             ^             4   2
  d       �     �   i        ���� � ������������i           ����             c             4   P
  �       �     �   i        ���� � ������������i           ����             h             5   n
  �       �	     �   i        ���� � ������������i           ����  
           V $           S   �
  �        �      �   j         ���� � ������������j           ����             [ (           U   "  f!       �     �   j         ���� � ������������j           ����             ` ,           W   ^  "       �     �   j         ���� � ������������j           ����             e 0           Y   �  �"       �     �   j        ���� � ������������j           ����             j 4           Z   �  �#       �     �   j        ���� � ������������j           ����             o 8           \     6$       �     �   j        ���� � ������������j           ����             t <           ^   N  �$       �     �   j        ���� � ������������j           ����             y @           `   �  �%       �     �   j        ���� � ������������j           ����             ~ D           b   �  R&       �     �   j        ���� � ������������j           ����             � H           c     '       �	     �   j        ���� � ������������j          ����             p 5          �   �  �7       �      �   k         ���� � ������������k          ����             u 9 !         �   L  09       �     �   k         ���� � ������������k          ����             z = $         �   �  �:       �     �   k         ���� � ������������k          ����              A '         �       <       �     �   k        ���� � ������������k          ����             � E *         �   Z  h=       �     �   k        ���� � ������������k          ����             � I -         �   �  �>       �     �   k        ���� � ������������k          ����             � M 0         �     8@       �     �   k        ���� � ������������k          ����             � Q 3         �   h  �A       �     �   k        ���� � ������������k          ����  ! "          � U 6         �   �  C       �     �   k        ���� � ������������k          ����  # $          � Y 9         �     pD       �	     �   k        ���� � ������������k          ����             � E &        �   �  �\       �      �   l         ���� � ������������l          ����             � I )        �   �  �^       �     �   l         ���� � ������������l          ����             � M ,         �   t  Da       �     �   l         ���� � ������������l          ����             � Q / #       �   �  �c       �     �   l        ���� � ������������l          ����             � U 2 &         d  �e       �     �   l        ���� � ������������l          ����              � Y 5 )         �  Lh       �     �   l        ���� � ������������l          ����  ! "          � ] 8 ,         T  �j       �     �   l        ���� � ������������l          ����  # $          � a ; /         �  �l       �     �   l        ���� � ������������l          ����  & '          � e > 2         D  To       �     �   l        ���� � ������������l          ����  ( )          � i A 5       #  �  �q       �	     �   l        ���� � ������������l           ����             / 3 4         2   `	  �       �      �   m         ���� � ������������m           ����             1 6 9         0   ~	  �       �     �   m         ���� � ������������m           ����             3 9 >         1   �	  8       �     �   m         ���� � ������������m           ����  	 
          5 < C         1   �	  t       �     �   m        ���� � ������������m           ����             7 ? H         2   �	  �       �     �   m        ���� � ������������m           ����             9 B M         3   �	  �       �     �   m        ���� � ������������m           ����             ; E R         3   
  (       �     �   m        ���� � ������������m           ����             = H W         4   2
  d       �     �   m        ���� � ������������m           ����             ? K \         4   P
  �       �     �   m        ���� � ������������m           ����             A N a         5   n
  �       �	     �   m        ���� � ������������m           ����             . ; O        S   �
  �        �      �   n         ���� � ������������n           ����  	 
          1 > T        U   "  f!       �     �   n         ���� � ������������n           ����             4 A Y        W   ^  "       �     �   n         ���� � ������������n           ����             7 D ^        Y   �  �"       �     �   n        ���� � ������������n           ����             : G c        Z   �  �#       �     �   n        ���� � ������������n           ����             = J h        \     6$       �     �   n        ���� � ������������n           ����             @ M m         ^   N  �$       �     �   n        ���� � ������������n           ����             C P r "       `   �  �%       �     �   n        ���� � ������������n           ����             F S w $       b   �  R&       �     �   n        ���� � ������������n           ����             I V | &       c     '       �	     �   n        ���� � ������������n          ����             6 B i        �   �  �7       �      �   o         ���� � ������������o          ����             9 F n        �   L  09       �     �   o         ���� � ������������o          ����             < J s        �   �  �:       �     �   o         ���� � ������������o          ����             ? N x !       �       <       �     �   o        ���� � ������������o          ����             B R } $       �   Z  h=       �     �   o        ���� � ������������o          ����             E V � '       �   �  �>       �     �   o        ���� � ������������o          ����             H Z � *       �     8@       �     �   o        ���� � ������������o          ����             K ^ � -       �   h  �A       �     �   o        ���� � ������������o          ����             N b � 0       �   �  C       �     �   o        ���� � ������������o          ����             Q f � 3       �     pD       �	     �   o        ���� � ������������o          ����             > S �         �   �  �\       �      �   p         ���� � ������������p          ����             A W � #       �   �  �^       �     �   p         ���� � ������������p          ����             D [ � &       �   t  Da       �     �   p         ���� � ������������p          ����             G _ � )       �   �  �c       �     �   p        ���� � ������������p          ����             J c � ,         d  �e       �     �   p        ���� � ������������p          ����             M g � /         �  Lh       �     �   p        ���� � ������������p          ����             P k � 2         T  �j       �     �   p        ���� � ������������p          ����             S o � 5         �  �l       �     �   p        ���� � ������������p          ����    !          V s � 8         D  To       �     �   p        ���� � ������������p          ����  " #          Y w � ;       #  �  �q       �	     �   p        ���� � ������������p           ����	              $             ����  .J       �      �� ��q         ���� � ������������q           ����	              )             ����.  \       �     �� ��q         ���� � ������������q           ����	              .             ����L  �       �     �� ��q         ���� � ������������q           ����	  
            3             ����j  �       �     �� ��q        ���� � ������������q           ����	              8             �����         �     �� ��q        ���� � ������������q           ����	              =             �����  L       �     �� ��q        ���� � ������������q           ����	              B             �����  �       �     �� ��q        ���� � ������������q           ����	              G             �����  �       �     �� ��q        ���� � ������������q           ����	              L             ����           �     �� ��q        ���� � ������������q           ����	              Q             ����  <       �	     �� ��q        ���� � ������������q           ����	   	           ? $           �����  �.       �      �� ��r         ���� � ������������r           ����	  
            D (           �����  v/       �     �� ��r         ���� � ������������r           ����	              I ,           ����  *0       �     �� ��r         ���� � ������������r           ����	              N 0           ����J  �0       �     �� ��r        ���� � ������������r           ����	              S 4           �����  �1       �     �� ��r        ���� � ������������r           ����	              X 8           �����  F2       �     �� ��r        ���� � ������������r           ����	              ] <           �����  �2       �     �� ��r        ���� � ������������r           ����	              b @           ����:  �3       �     �� ��r        ���� � ������������r           ����	              g D           ����v  b4       �     �� ��r        ���� � ������������r           ����	              l H           �����  5       �	     �� ��r        ���� � ������������r          ����	              Y 5          �����  �J       �      �� ��s         ���� � ������������s          ����	              ^ 9 !         �����  �K       �     �� ��s         ���� � ������������s          ����	              c = $         ����V  XM       �     �� ��s         ���� � ������������s          ����	              h A '         �����  �N       �     �� ��s        ���� � ������������s          ����	              m E *         ����
  (P       �     �� ��s        ���� � ������������s          ����	              r I -         ����d  �Q       �     �� ��s        ���� � ������������s          ����	              w M 0         �����  �R       �     �� ��s        ���� � ������������s          ����	              | Q 3         ����  `T       �     �� ��s        ���� � ������������s          ����	               � U 6         ����r  �U       �     �� ��s        ���� � ������������s          ����	  ! "           � Y 9         �����  0W       �	     �� ��s        ���� � ������������s          ����	              r E &        ����4  t       �      �� ��t         ���� � ������������t          ����	              x I )        �����  \v       �     �� ��t         ���� � ������������t          ����	              ~ M ,         ����$  �x       �     �� ��t         ���� � ������������t          ����	              � Q / #       �����  {       �     �� ��t        ���� � ������������t          ����	              � U 2 &       ����  d}       �     �� ��t        ���� � ������������t          ����	              � Y 5 )       �����  �       �     �� ��t        ���� � ������������t          ����	               � ] 8 ,       ����  �       �     �� ��t        ���� � ������������t          ����	  ! "           � a ; /       ����|  l�       �     �� ��t        ���� � ������������t          ����	  $ %           � e > 2       �����  Ć       �     �� ��t        ���� � ������������t          ����	  & '           � i A 5       ����l  �       �	     �� ��t        ���� � ������������t           ����	                         ����  .J       �      �� ��u         ���� � ������������u           ����	                "         ����.  \       �     �� ��u         ���� � ������������u           ����	               " '         ����L  �       �     �� ��u         ���� � ������������u           ����	   	            % ,         ����j  �       �     �� ��u        ���� � ������������u           ����	  
            ! ( 1         �����         �     �� ��u        ���� � ������������u           ����	              # + 6         �����  L       �     �� ��u        ���� � ������������u           ����	              % . ;         �����  �       �     �� ��u        ���� � ������������u           ����	              ' 1 @         �����  �       �     �� ��u        ���� � ������������u           ����	              ) 4 E         ����           �     �� ��u        ���� � ������������u           ����	              + 7 J         ����  <       �	     �� ��u        ���� � ������������u           ����	               $ 8        �����  �.       �      �� ��v         ���� � ������������v           ����	   	            ' =        �����  v/       �     �� ��v         ���� � ������������v           ����	  
             * B        ����  *0       �     �� ��v         ���� � ������������v           ����	              ! - G        ����J  �0       �     �� ��v        ���� � ������������v           ����	              $ 0 L        �����  �1       �     �� ��v        ���� � ������������v           ����	              ' 3 Q        �����  F2       �     �� ��v        ���� � ������������v           ����	              * 6 V         �����  �2       �     �� ��v        ���� � ������������v           ����	              - 9 [ "       ����:  �3       �     �� ��v        ���� � ������������v           ����	              0 < ` $       ����v  b4       �     �� ��v        ���� � ������������v           ����	              3 ? e &       �����  5       �	     �� ��v        ���� � ������������v          ����	  
              + R        �����  �J       �      �� ��w         ���� � ������������w          ����	              # / W        �����  �K       �     �� ��w         ���� � ������������w          ����	              & 3 \        ����V  XM       �     �� ��w         ���� � ������������w          ����	              ) 7 a !       �����  �N       �     �� ��w        ���� � ������������w          ����	              , ; f $       ����
  (P       �     �� ��w        ���� � ������������w          ����	              / ? k '       ����d  �Q       �     �� ��w        ���� � ������������w          ����	              2 C p *       �����  �R       �     �� ��w        ���� � ������������w          ����	              5 G u -       ����  `T       �     �� ��w        ���� � ������������w          ����	              8 K z 0       ����r  �U       �     �� ��w        ���� � ������������w          ����	              ; O  3       �����  0W       �	     �� ��w        ���� � ������������w          ����	              ( < k         ����4  t       �      �� ��x         ���� � ������������x          ����	              + @ q #       �����  \v       �     �� ��x         ���� � ������������x          ����	              . D w &       ����$  �x       �     �� ��x         ���� � ������������x          ����	              1 H } )       �����  {       �     �� ��x        ���� � ������������x          ����	              4 L � ,       ����  d}       �     �� ��x        ���� � ������������x          ����	              7 P � /       �����  �       �     �� ��x        ���� � ������������x          ����	              : T � 2       ����  �       �     �� ��x        ���� � ������������x          ����	              = X � 5       ����|  l�       �     �� ��x        ���� � ������������x          ����	               @ \ � 8       �����  Ć       �     �� ��x        ���� � ������������x          ����	  ! "           C ` � ;       ����l  �       �	     �� ��x        ���� � ������������x           ����
              1             �����  t1       7      �� ��y         ���� � ������������y           ����
              6             �����  <       7     �� ��y         ���� � ������������y           ����
   	           ;             �����  x       7     �� ��y         ���� � ������������y           ����
              @             �����  �       7     �� ��y        ���� � ������������y           ����
              E             �����  �       7     �� ��y        ���� � ������������y           ����
              J             ����  ,       7     �� ��y        ���� � ������������y           ����
              O             ����4  h       7     �� ��y        ���� � ������������y           ����
              T             ����R  �       7     �� ��y        ���� � ������������y           ����
              Y             ����p  �       7     �� ��y        ���� � ������������y           ����
              ^             �����         7	     �� ��y        ���� � ������������y           ����
  	 
           L $           ����  *       8      �� ��z         ���� � ������������z           ����
              Q (           ����B  �*       8     �� ��z         ���� � ������������z           ����
              V ,           ����~  z+       8     �� ��z         ���� � ������������z           ����
              [ 0           �����  .,       8     �� ��z        ���� � ������������z           ����
              ` 4           �����  �,       8     �� ��z        ���� � ������������z           ����
              e 8           ����2  �-       8     �� ��z        ���� � ������������z           ����
              j <           ����n  J.       8     �� ��z        ���� � ������������z           ����
              o @           �����  �.       8     �� ��z        ���� � ������������z           ����
              t D           �����  �/       8     �� ��z        ���� � ������������z           ����
              y H           ����"  f0       8	     �� ��z        ���� � ������������z          ����
              f 5          ����  HD       9      �� ��{         ���� � ������������{          ����
              k 9 !         ����l  �E       9     �� ��{         ���� � ������������{          ����
              p = $         �����  G       9     �� ��{         ���� � ������������{          ����
              u A '         ����   �H       9     �� ��{        ���� � ������������{          ����
              z E *         ����z  �I       9     �� ��{        ���� � ������������{          ����
               I -         �����  PK       9     �� ��{        ���� � ������������{          ����
              � M 0         ����.  �L       9     �� ��{        ���� � ������������{          ����
              � Q 3         �����   N       9     �� ��{        ���� � ������������{          ����
    !           � U 6         �����  �O       9     �� ��{        ���� � ������������{          ����
  " #           � Y 9         ����<  �P       9	     �� ��{        ���� � ������������{          ����
               E &        �����  4l       :      �� ��|         ���� � ������������|          ����
              � I )        ����  �n       :     �� ��|         ���� � ������������|          ����
              � M ,         �����  �p       :     �� ��|         ���� � ������������|          ����
              � Q / #       ����  <s       :     �� ��|        ���� � ������������|          ����
              � U 2 &       �����  �u       :     �� ��|        ���� � ������������|          ����
              � Y 5 )       �����  �w       :     �� ��|        ���� � ������������|          ����
    !           � ] 8 ,       ����t  Dz       :     �� ��|        ���� � ������������|          ����
  " #           � a ; /       �����  �|       :     �� ��|        ���� � ������������|          ����
  % &           � e > 2       ����d  �~       :     �� ��|        ���� � ������������|          ����
  ' (           � i A 5       �����  L�       :	     �� ��|        ���� � ������������|           ����
              & ) *         �����  t1       F      �� ��}         ���� � ������������}           ����
              ( , /         �����  <       F     �� ��}         ���� � ������������}           ����
              * / 4         �����  x       F     �� ��}         ���� � ������������}           ����
   	           , 2 9         �����  �       F     �� ��}        ���� � ������������}           ����
  
            . 5 >         �����  �       F     �� ��}        ���� � ������������}           ����
              0 8 C         ����  ,       F     �� ��}        ���� � ������������}           ����
              2 ; H         ����4  h       F     �� ��}        ���� � ������������}           ����
              4 > M         ����R  �       F     �� ��}        ���� � ������������}           ����
              6 A R         ����p  �       F     �� ��}        ���� � ������������}           ����
              8 D W         �����         F	     �� ��}        ���� � ������������}           ����
              % 1 E        ����  *       G      �� ��~         ���� � ������������~           ����
   	           ( 4 J        ����B  �*       G     �� ��~         ���� � ������������~           ����
  
            + 7 O        ����~  z+       G     �� ��~         ���� � ������������~           ����
              . : T        �����  .,       G     �� ��~        ���� � ������������~           ����
              1 = Y        �����  �,       G     �� ��~        ���� � ������������~           ����
              4 @ ^        ����2  �-       G     �� ��~        ���� � ������������~           ����
              7 C c         ����n  J.       G     �� ��~        ���� � ������������~           ����
              : F h "       �����  �.       G     �� ��~        ���� � ������������~           ����
              = I m $       �����  �/       G     �� ��~        ���� � ������������~           ����
              @ L r &       ����"  f0       G	     �� ��~        ���� � ������������~          ����
  
            - 8 _        ����  HD       H      �� ��         ���� � ������������          ����
              0 < d        ����l  �E       H     �� ��         ���� � ������������          ����
              3 @ i        �����  G       H     �� ��         ���� � ������������          ����
              6 D n !       ����   �H       H     �� ��        ���� � ������������          ����
              9 H s $       ����z  �I       H     �� ��        ���� � ������������          ����
              < L x '       �����  PK       H     �� ��        ���� � ������������          ����
              ? P } *       ����.  �L       H     �� ��        ���� � ������������          ����
              B T � -       �����   N       H     �� ��        ���� � ������������          ����
              E X � 0       �����  �O       H     �� ��        ���� � ������������          ����
              H \ � 3       ����<  �P       H	     �� ��        ���� � ������������          ����
              5 I x         �����  4l       I      �� ���         ���� � �������������          ����
              8 M ~ #       ����  �n       I     �� ���         ���� � �������������          ����
              ; Q � &       �����  �p       I     �� ���         ���� � �������������          ����
              > U � )       ����  <s       I     �� ���        ���� � �������������          ����
              A Y � ,       �����  �u       I     �� ���        ���� � �������������          ����
              D ] � /       �����  �w       I     �� ���        ���� � �������������          ����
              G a � 2       ����t  Dz       I     �� ���        ���� � �������������          ����
              J e � 5       �����  �|       I     �� ���        ���� � �������������          ����
               M i � 8       ����d  �~       I     �� ���        ���� � �������������          ����
  ! "           P m � ;       �����  L�       I	     �� ���        ���� � �������������           ����              >             �����  X       �      �� ���         ���� � �������������           ����              C             ����  $       �     �� ���         ���� � �������������           ����  	 
           H             ����0  `       �     �� ���         ���� � �������������           ����              M             ����N  �       �     �� ���        ���� � �������������           ����              R             ����l  �       �     �� ���        ���� � �������������           ����              W             �����         �     �� ���        ���� � �������������           ����              \             �����  P       �     �� ���        ���� � �������������           ����              a             �����  �       �     �� ���        ���� � �������������           ����              f             �����  �       �     �� ���        ���� � �������������           ����              k             ����         �	     �� ���        ���� � �������������           ����  
            Y $           ����z  n
       �      �� ���         ���� � �������������           ����              ^ (           �����  "       �     �� ���         ���� � �������������           ����              c ,           �����  �       �     �� ���         ���� � �������������           ����              h 0           ����.  �       �     �� ���        ���� � �������������           ����              m 4           ����j  >       �     �� ���        ���� � �������������           ����              r 8           �����  �       �     �� ���        ���� � �������������           ����              w <           �����  �       �     �� ���        ���� � �������������           ����              | @           ����  Z       �     �� ���        ���� � �������������           ����              � D           ����Z         �     �� ���        ���� � �������������           ����              � H           �����  �       �	     �� ���        ���� � �������������          ����              s 5          �����         �      �� ���         ���� � �������������          ����              x 9 !         �����  �       �     �� ���         ���� � �������������          ����              } = $         ����:  �       �     �� ���         ���� � �������������          ����              � A '         �����  P       �     �� ���        ���� � �������������          ����              � E *         �����  �       �     �� ���        ���� � �������������          ����              � I -         ����H   !       �     �� ���        ���� � �������������          ����              � M 0         �����  �"       �     �� ���        ���� � �������������          ����              � Q 3         �����  �#       �     �� ���        ���� � �������������          ����  ! "           � U 6         ����V	  X%       �     �� ���        ���� � �������������          ����  # $           � Y 9         �����	  �&       �	     �� ���        ���� � �������������          ����              � E &        ����  x7       �      �� ���         ���� � �������������          ����              � I )        �����  �9       �     �� ���         ���� � �������������          ����              � M ,         ����  (<       �     �� ���         ���� � �������������          ����              � Q / #       �����  �>       �     �� ���        ���� � �������������          ����              � U 2 &       �����  �@       �     �� ���        ���� � �������������          ����               � Y 5 )       ����p  0C       �     �� ���        ���� � �������������          ����  ! "           � ] 8 ,       �����  �E       �     �� ���        ���� � �������������          ����  # $           � a ; /       ����`  �G       �     �� ���        ���� � �������������          ����  & '           � e > 2       �����  8J       �     �� ���        ���� � �������������          ����  ( )           � i A 5       ����P  �L       �	     �� ���        ���� � �������������           ����              2 6 7         �����  X       �      �� ���         ���� � �������������           ����              4 9 <         ����  $       �     �� ���         ���� � �������������           ����              6 < A         ����0  `       �     �� ���         ���� � �������������           ����  	 
           8 ? F         ����N  �       �     �� ���        ���� � �������������           ����              : B K         ����l  �       �     �� ���        ���� � �������������           ����              < E P         �����         �     �� ���        ���� � �������������           ����              > H U         �����  P       �     �� ���        ���� � �������������           ����              @ K Z         �����  �       �     �� ���        ���� � �������������           ����              B N _         �����  �       �     �� ���        ���� � �������������           ����              D Q d         ����         �	     �� ���        ���� � �������������           ����              1 > R        ����z  n
       �      �� ���         ���� � �������������           ����  	 
           4 A W        �����  "       �     �� ���         ���� � �������������           ����              7 D \        �����  �       �     �� ���         ���� � �������������           ����              : G a        ����.  �       �     �� ���        ���� � �������������           ����              = J f        ����j  >       �     �� ���        ���� � �������������           ����              @ M k        �����  �       �     �� ���        ���� � �������������           ����              C P p         �����  �       �     �� ���        ���� � �������������           ����              F S u "       ����  Z       �     �� ���        ���� � �������������           ����              I V z $       ����Z         �     �� ���        ���� � �������������           ����              L Y  &       �����  �       �	     �� ���        ���� � �������������          ����              9 E l        �����         �      �� ���         ���� � �������������          ����              < I q        �����  �       �     �� ���         ���� � �������������          ����              ? M v        ����:  �       �     �� ���         ���� � �������������          ����              B Q { !       �����  P       �     �� ���        ���� � �������������          ����              E U � $       �����  �       �     �� ���        ���� � �������������          ����              H Y � '       ����H   !       �     �� ���        ���� � �������������          ����              K ] � *       �����  �"       �     �� ���        ���� � �������������          ����              N a � -       �����  �#       �     �� ���        ���� � �������������          ����              Q e � 0       ����V	  X%       �     �� ���        ���� � �������������          ����              T i � 3       �����	  �&       �	     �� ���        ���� � �������������          ����              A V �         ����  x7       �      �� ���         ���� � �������������          ����              D Z � #       �����  �9       �     �� ���         ���� � �������������          ����              G ^ � &       ����  (<       �     �� ���         ���� � �������������          ����              J b � )       �����  �>       �     �� ���        ���� � �������������          ����              M f � ,       �����  �@       �     �� ���        ���� � �������������          ����              P j � /       ����p  0C       �     �� ���        ���� � �������������          ����              S n � 2       �����  �E       �     �� ���        ���� � �������������          ����              V r � 5       ����`  �G       �     �� ���        ���� � �������������          ����    !           Y v � 8       �����  8J       �     �� ���        ���� � �������������          ����  " #           \ z � ;       ����P  �L       �	     �� ���        ���� � �������������           ����              K             �����  �        �      �� ���         ���� � �������������           ����   	           P             �����  |       �     �� ���         ���� � �������������           ����  
            U             �����  �       �     �� ���         ���� � �������������           ����              Z             �����  �       �     �� ���        ���� � �������������           ����              _             ����  0        �     �� ���        ���� � �������������           ����              d             ����6  l        �     �� ���        ���� � �������������           ����              i             ����T  �        �     �� ���        ���� � �������������           ����              n             ����r  �        �     �� ���        ���� � �������������           ����              s             �����   !       �     �� ���        ���� � �������������           ����              x             �����  \!       �	     �� ���        ���� � �������������           ����              f $           ����&  r3       �      �� ���         ���� � �������������           ����              k (           ����b  &4       �     �� ���         ���� � �������������           ����              p ,           �����  �4       �     �� ���         ���� � �������������           ����              u 0           �����  �5       �     �� ���        ���� � �������������           ����              z 4           ����  B6       �     �� ���        ���� � �������������           ����               8           ����R  �6       �     �� ���        ���� � �������������           ����              � <           �����  �7       �     �� ���        ���� � �������������           ����              � @           �����  ^8       �     �� ���        ���� � �������������           ����              � D           ����  9       �     �� ���        ���� � �������������           ����               � H           ����B  �9       �	     �� ���        ���� � �������������          ����              � 5          ����2  �P       �      �� ���         ���� � �������������          ����              � 9 !         �����  0R       �     �� ���         ���� � �������������          ����              � = $         �����  �S       �     �� ���         ���� � �������������          ����              � A '         ����@   U       �     �� ���        ���� � �������������          ����              � E *         �����  hV       �     �� ���        ���� � �������������          ����              � I -         �����  �W       �     �� ���        ���� � �������������          ����              � M 0         ����N  8Y       �     �� ���        ���� � �������������          ����               � Q 3         �����  �Z       �     �� ���        ���� � �������������          ����  " #           � U 6         ����  \       �     �� ���        ���� � �������������          ����  $ %           � Y 9         ����\  p]       �	     �� ���        ���� � �������������          ����              � E &        �����  �{       �      �� ���         ���� � �������������          ����              � I )        ����<  ,~       �     �� ���         ���� � �������������          ����              � M ,         �����  ��       �     �� ���         ���� � �������������          ����              � Q / #       ����,  ܂       �     �� ���        ���� � �������������          ����              � U 2 &       �����  4�       �     �� ���        ���� � �������������          ����    !           � Y 5 )       ����  ��       �     �� ���        ���� � �������������          ����  " #           � ] 8 ,       �����  �       �     �� ���        ���� � �������������          ����  $ %           � a ; /       ����  <�       �     �� ���        ���� � �������������          ����  ' (           � e > 2       �����  ��       �     �� ���        ���� � �������������          ����  ) *           � i A 5       �����  �       �	     �� ���        ���� � �������������           ����              ? C D         �����  �        �      �� ���         ���� � �������������           ����              A F I         �����  |       �     �� ���         ���� � �������������           ����              C I N         �����  �       �     �� ���         ���� � �������������           ����  	 
           E L S         �����  �       �     �� ���        ���� � �������������           ����              G O X         ����  0        �     �� ���        ���� � �������������           ����              I R ]         ����6  l        �     �� ���        ���� � �������������           ����              K U b         ����T  �        �     �� ���        ���� � �������������           ����              M X g         ����r  �        �     �� ���        ���� � �������������           ����              O [ l         �����   !       �     �� ���        ���� � �������������           ����              Q ^ q         �����  \!       �	     �� ���        ���� � �������������           ����              > K _        ����&  r3       �      �� ���         ���� � �������������           ����  	 
           A N d        ����b  &4       �     �� ���         ���� � �������������           ����              D Q i        �����  �4       �     �� ���         ���� � �������������           ����              G T n        �����  �5       �     �� ���        ���� � �������������           ����              J W s        ����  B6       �     �� ���        ���� � �������������           ����              M Z x        ����R  �6       �     �� ���        ���� � �������������           ����              P ] }         �����  �7       �     �� ���        ���� � �������������           ����              S ` � "       �����  ^8       �     �� ���        ���� � �������������           ����              V c � $       ����  9       �     �� ���        ���� � �������������           ����              Y f � &       ����B  �9       �	     �� ���        ���� � �������������          ����              F R y        ����2  �P       �      �� ���         ���� � �������������          ����              I V ~        �����  0R       �     �� ���         ���� � �������������          ����              L Z �        �����  �S       �     �� ���         ���� � �������������          ����              O ^ � !       ����@   U       �     �� ���        ���� � �������������          ����              R b � $       �����  hV       �     �� ���        ���� � �������������          ����              U f � '       �����  �W       �     �� ���        ���� � �������������          ����              X j � *       ����N  8Y       �     �� ���        ���� � �������������          ����              [ n � -       �����  �Z       �     �� ���        ���� � �������������          ����              ^ r � 0       ����  \       �     �� ���        ���� � �������������          ����              a v � 3       ����\  p]       �	     �� ���        ���� � �������������          ����              N c �         �����  �{       �      �� ���         ���� � �������������          ����              Q g � #       ����<  ,~       �     �� ���         ���� � �������������          ����              T k � &       �����  ��       �     �� ���         ���� � �������������          ����              W o � )       ����,  ܂       �     �� ���        ���� � �������������          ����              Z s � ,       �����  4�       �     �� ���        ���� � �������������          ����              ] w � /       ����  ��       �     �� ���        ���� � �������������          ����              ` { � 2       �����  �       �     �� ���        ���� � �������������          ����              c  � 5       ����  <�       �     �� ���        ���� � �������������          ����    !           f � � 8       �����  ��       �     �� ���        ���� � �������������          ����  " #           i � � ;       �����  �       �	     �� ���        ���� � �������������           ����              N             ����0  �        E      �� ���         ���� � �������������           ����   	           S             ����N  �"       E     �� ���         ���� � �������������           ����  
            X             ����l  �"       E     �� ���         ���� � �������������           ����              ]             �����  #       E     �� ���        ���� � �������������           ����              b             �����  P#       E     �� ���        ���� � �������������           ����              g             �����  �#       E     �� ���        ���� � �������������           ����              l             �����  �#       E     �� ���        ���� � �������������           ����              q             ����  $       E     �� ���        ���� � �������������           ����              v             ����   @$       E     �� ���        ���� � �������������           ����              {             ����>  |$       E	     �� ���        ���� � �������������           ����              i $           �����  "8       F      �� ���         ���� � �������������           ����              n (           �����  �8       F     �� ���         ���� � �������������           ����              s ,           ����.  �9       F     �� ���         ���� � �������������           ����              x 0           ����j  >:       F     �� ���        ���� � �������������           ����              } 4           �����  �:       F     �� ���        ���� � �������������           ����              � 8           �����  �;       F     �� ���        ���� � �������������           ����              � <           ����  Z<       F     �� ���        ���� � �������������           ����              � @           ����Z  =       F     �� ���        ���� � �������������           ����              � D           �����  �=       F     �� ���        ���� � �������������           ����               � H           �����  v>       F	     �� ���        ���� � �������������          ����              � 5          �����  W       G      �� ���         ���� � �������������          ����              � 9 !         ����  pX       G     �� ���         ���� � �������������          ����              � = $         ����v  �Y       G     �� ���         ���� � �������������          ����              � A '         �����  @[       G     �� ���        ���� � �������������          ����              � E *         ����*  �\       G     �� ���        ���� � �������������          ����              � I -         �����  ^       G     �� ���        ���� � �������������          ����              � M 0         �����  x_       G     �� ���        ���� � �������������          ����               � Q 3         ����8  �`       G     �� ���        ���� � �������������          ����  " #           � U 6         �����  Hb       G     �� ���        ���� � �������������          ����  $ %           � Y 9         �����  �c       G	     �� ���        ���� � �������������          ����              � E &        ����T  ��       H      �� ���         ���� � �������������          ����              � I )        �����  ��       H     �� ���         ���� � �������������          ����              � M ,         ����D  T�       H     �� ���         ���� � �������������          ����              � Q / #       �����  ��       H     �� ���        ���� � �������������          ����              � U 2 &       ����4  �       H     �� ���        ���� � �������������          ����    !           � Y 5 )       �����  \�       H     �� ���        ���� � �������������          ����  " #           � ] 8 ,       ����$  ��       H     �� ���        ���� � �������������          ����  $ %           � a ; /       �����  �       H     �� ���        ���� � �������������          ����  ' (           � e > 2       ����  d�       H     �� ���        ���� � �������������          ����  ) *           � i A 5       �����  ��       H	     �� ���        ���� � �������������           ����              B F G         ����0  �        T      �� ���         ���� � �������������           ����              D I L         ����N  �"       T     �� ���         ���� � �������������           ����              F L Q         ����l  �"       T     �� ���         ���� � �������������           ����  	 
           H O V         �����  #       T     �� ���        ���� � �������������           ����              J R [         �����  P#       T     �� ���        ���� � �������������           ����              L U `         �����  �#       T     �� ���        ���� � �������������           ����              N X e         �����  �#       T     �� ���        ���� � �������������           ����              P [ j         ����  $       T     �� ���        ���� � �������������           ����              R ^ o         ����   @$       T     �� ���        ���� � �������������           ����              T a t         ����>  |$       T	     �� ���        ���� � �������������           ����              A N b        �����  "8       U      �� ���         ���� � �������������           ����  	 
           D Q g        �����  �8       U     �� ���         ���� � �������������           ����              G T l        ����.  �9       U     �� ���         ���� � �������������           ����              J W q        ����j  >:       U     �� ���        ���� � �������������           ����              M Z v        �����  �:       U     �� ���        ���� � �������������           ����              P ] {        �����  �;       U     �� ���        ���� � �������������           ����              S ` �         ����  Z<       U     �� ���        ���� � �������������           ����              V c � "       ����Z  =       U     �� ���        ���� � �������������           ����              Y f � $       �����  �=       U     �� ���        ���� � �������������           ����              \ i � &       �����  v>       U	     �� ���        ���� � �������������          ����              I U |        �����  W       V      �� ���         ���� � �������������          ����              L Y �        ����  pX       V     �� ���         ���� � �������������          ����              O ] �        ����v  �Y       V     �� ���         ���� � �������������          ����              R a � !       �����  @[       V     �� ���        ���� � �������������          ����              U e � $       ����*  �\       V     �� ���        ���� � �������������          ����              X i � '       �����  ^       V     �� ���        ���� � �������������          ����              [ m � *       �����  x_       V     �� ���        ���� � �������������          ����              ^ q � -       ����8  �`       V     �� ���        ���� � �������������          ����              a u � 0       �����  Hb       V     �� ���        ���� � �������������          ����              d y � 3       �����  �c       V	     �� ���        ���� � �������������          ����              Q f �         ����T  ��       W      �� ���         ���� � �������������          ����              T j � #       �����  ��       W     �� ���         ���� � �������������          ����              W n � &       ����D  T�       W     �� ���         ���� � �������������          ����              Z r � )       �����  ��       W     �� ���        ���� � �������������          ����              ] v � ,       ����4  �       W     �� ���        ���� � �������������          ����              ` z � /       �����  \�       W     �� ���        ���� � �������������          ����              c ~ � 2       ����$  ��       W     �� ���        ���� � �������������          ����              f � � 5       �����  �       W     �� ���        ���� � �������������          ����    !           i � � 8       ����  d�       W     �� ���        ���� � �������������          ����  " #           l � � ;       �����  ��       W	     �� ���        ���� � �������������            ��d ���                          �      ]         �  
   ��, ���         ������  ����������������         ��d ���                         �   <   �         �  
   ��, ���         ������  ����������������         ��d ���                         �   _           �  
   ��, ���         ������  ����������������         ��d ��L                         �   �   �        �  
   ��, ���         ������  ����������������         ��e ���                          �   %   q         �     ��- ���         ������  ����������������         ��e ���                         �   >   �         �     ��- ���         ������  ����������������         ��e ���                         �   _           �     ��- ���         ������  ����������������         ��e ��L                         �   �   �        �     ��- ���         ������  ����������������         ��f ��-                          �   (   }         �      ��, ���         ������  ����������������         ��f ��7                          �   ?   �         �      ��, ���         ������  ����������������         ��f ��A                          �   `            �      ��, ���         ������  ����������������         ��f ��K                          �   �   �        �      ��, ���         ������  ����������������          g                             �����   �        �      ��$ ���         ����   ����������������         g                            ����B  �        �      ��$ ���         ����   ����������������         g                            ����[  l        �      ��$ ���         ����   ����������������         g                +          ����'  �#        �      ��$ ���         ����   ����������������         g                D "         �����
  �?        �      ��$ ���         ����   ����������������         g                O 1 & "       �����  �g        �      ��$ ���         ����   ����������������         g                [ @ . )       �����  �        �      ��$ ���         ����   ����������������         g                h Q 7 1       ����U  ��        �      ��$ ���         ����   ����������������         g                x c A :       �����  @<       �      ��$ ���         ����	   ����������������        	 g                � | L A       �����&  ʨ       �      ��$ ���         ����
   ����������������        
 g                � � X L       ����O.  �+       �      ��$ ���         ����   ����������������         g                � � e U       �����6  �       �      ��$ ���         ����   ����������������         g                           �����   �        �      ��% ���         ����   ����������������         g                          ����B  �        �      ��% ���         ����   ����������������         g                  %        ����[  l        �      ��% ���         ����   ����������������         g                  4        ����'  �#        �      ��% ���         ����   ����������������         g                " % >        �����
  �?        �      ��% ���         ����   ����������������         g                1 6 U "       �����  �g        �      ��% ���         ����   ����������������         g                @ @ b )       �����  �        �      ��% ���         ����   ����������������         g                Q W  1       ����U  ��        �      ��% ���         ����   ����������������         g                c d � :       �����  @<       �      ��% ���         ����	   ����������������          g                v � � A       �����&  ʨ       �      ��% ���         ����
   ����������������        ! g                � � � L       ����O.  �+       �      ��% ���         ����   ����������������        " g                � � � U       �����6  �       �      ��% ���         ����   ����������������       ����� ��                            �����   �        T      ��7 ���         ������  ����������������       ����� ��                           ����B  �        U      ��7 ���         ������  ����������������       ����� ��                           ����[  l        V      ��7 ���         ������  ����������������       ����� ��                           ����'  �#        W      ��7 ���         ������  ����������������       ����� ��                           �����
  �?        X      ��7 ���         ������  ����������������       ����� ��                           �����  x        Y      ��8 ���         ������  ����������������       ����� ��                           ����  Z	        Z      ��8 ���         ������  ����������������       ����� ��                           ����7  �        [      ��8 ���         ������  ����������������       ����� ��                           ����  (        \      ��8 ���         ������  ����������������       ����� ��            	               �����  E        ]      ��8 ���         ������  ����������������       ����� ��            
               �����  4        ^      ��9 ���         ������  ����������������       ����� ��                           �����  �        _      ��9 ���         ������  ����������������       ����� ��                           ����  L        `      ��9 ���         ������  ����������������       ����� ��                           �����  [,        a      ��9 ���         ������  ����������������       ����� ��                           ����^  4J        b      ��9 ���         ������  ����������������        ����� ��                            ����                   ��> ���         ������  ����������������           ��@Iv2    � � J >         �,  |�                 �     +..���� � �����  �  �              ��LV�2    � � N B         �-  �                �     +..���� � �����  �  �              ��+Xc�2    � � R F       /  |.  \�                �     +..���� � �����  �  �              ��7dp�2    � � V J       D  l/  ̪                �    +..���� � �����  �  �              ��Cp}�2    � � Z N       Z  \0  <�                �    +..���� � �����  �  �              ��O|��2     � ^ R       o  L1  ��                �    +..���� � �����  �  �              ��[���2    � b V       �  <2  �                �    +..���� � �����  �  �              ��g���2    � f Z       �  ,3  ��                �    +..���� � �����  �  �              ��s���2    � j ^       �  4  ��                �    +..���� � �����  �  �              �����2    � n b       �  5  l�   
    	         �    +..���� � �����  �  �             ��]���2    � Y M       �  �8  �7      	           �     G������	 � �����  �  �             ��j���2    � ] Q       �  �9  �B      	          �     G������	 � �����  �  �             ��w���2    � a U       �  �:  M      	          �     G������	 � �����  �  �             �����2    � e Y       �  �;  �W      	          �    G������	 � �����  �  �             �����2    � i ]         =  (b      	          �    G������	 � �����  �  �             �����'2    $� m a       5  >  �l      	          �    G������	 � �����  �  �             �����72    +� q e       P   ?  @w      	          �    G������	 � �����  �  �             ����G2    2� u i       k  .@  ́      	          �    G������	 � �����  �  �             ����W2    9� y m       �  <A  X�   	   	          �    G������	 � �����  �  �             ���$g2    @� } q       �  JB  �      	 	         �    G������	 � �����  �  �             ���� G2    )� h \       �  �F  �      
       	    �     �������
 � �����  �  �             ����X2    0� l `       �  �G  z      
      	    �     �������
 � �����  �  �             ���"i2    7� p d         �H  ^!      
      	    �     �������
 � �����  �  �             ���3z2    >� t h       $  J  B.      
      	    �    �������
 � �����  �  �             ���%D�2    E� x l       E  2K  &;      
      	    �    �������
 � �����  �  �             ���4U�2    L� | p       f  ^L  
H      
      	    �    �������
 � �����  �  �             ��Cf�2    S� � t       �  �M  �T   
   
      	    �    �������
 � �����  �  �             ��Rw�2    Z� � x       �  �N  �a   	   
      	    �    �������
 � �����  �  �             ��$a��2    a� � |       �  �O  �n      
      	    �    �������
 � �����  �  �             ��3p��2    h� � �       �  Q  �{      
 	     	    �    �������
 � �����  �  �             ��	Iq�2    P� v j       J
  �U  �             
    �     ɖ����� � �����  �  �             ��Z��2    W� { o       q
  W  `            
    �     ɖ����� � �����  �  �             ��)k��2    ^� � t       �
  RX  �#            
    �     ɖ����� � �����  �  �             ��9|��2    e� � y       �
  �Y  P3            
    �    ɖ����� � �����  �  �             ��I��2    l� � ~       �
  �Z  �B            
    �    ɖ����� � �����  �  �             ��Y��2    s� � �         0\  @R   	         
    �    ɖ����� � �����  �  �             ��i��-2    z � �       7  z]  �a            
    �    ɖ����� � �����  �  �             ��y��@2    �� �       _  �^  0q            
    �    ɖ����� � �����  �  �             ����S2    �� �       �  `  ��            
    �    ɖ����� � �����  �  �             ����f2    �� �       �  Xa   �       	     
    �    ɖ����� � �����  �  �             ��j��>2    v� � �       S  �f  �4                 �     �m����� � �����  �  �             ��{��S2    } � �       �  �g  �F                �     �m����� � �����  �  �             ����h2    �� �       �  Pi  Y                �     �m����� � �����  �  �             ����"}2    �� �       �  �j  Xk   
             �    �m����� � �����  �  �             ��� 6�2    �� �          l  �}   	             �    �m����� � �����  �  �             ���J�2    �� �       =  �m  �                �    �m����� � �����  �  �             ���$^�2    �� �       l  �n  0�                �    �m����� � �����  �  �             ���6r�2    �$� �       �  Xp  x�                �    �m����� � �����  �  �             ���H��2    �*� �       �  �q  ��                �    �m����� � �����  �  �             ��Z��2    �0� �       �  (s  �       	         �    �m����� �    �  �  �             ���+i�2    �� �       �  �x  �                 �     TX����� � �����  �  �             ���?~�2    �� �         Nz  D�                �     TX����� � �����  �  �             ���S��2    �#� �       V  �{  ��   	             �     TX����� � �����  �  �             ��g�2    �)� �       �  Z}  ��                �    TX����� � �����  �  �             ��{�'2    �/� �       �  �~  @�                �    TX����� � �����  �  �             ��.��=2    �5� �       �  f�  �                �    TX����� � �����  �  �             ��A��S2    �;� �       0  �  �                �    TX����� � �����  �  �             ��T��i2    �A� �       g  r�  <0                �    TX����� � �����  �  �             ��g�2    �G� �       �  ��  �E                �    TX����� � �����  �  �             ��z�&�2    �M� �       �  ~�  �Z        	         �    TX����� �    �  �  �             ��C��e2    �4� �         ��  �<   
              �     :������ � �����  �  �             ��W�}2    �;� �       U  :�  fU   	             �     :������ � �����  �  �             ��k��2    �B� �       �  ޏ  n                �     :������ � �����  �  �             ���6�2    �I� �       �  ��  ��                �    :������ � �����  �  �             ���M�2    �P� �         &�  :�                �    :������ � �����  �  �             ���d�2    �W� �       Q  ʔ  ַ                �    :������ � �����  �  �             ���+{�2    �^� �       �  n�  r�                �    :������ � �����  �  �             ���@�2    e� �       �  �  �                �    :������ � �����  �  �             ���U�%2    
l� �         ��  �	   ��            �    :������ � �����  �  �             ���j�=2    s� �       M  Z�  F	   ��   	         �    :������ �    �  �  �             ���3�	2    �Z� �       �  �  �
                 �     �Z���� � �����  �  �             ���J�#2     a� �       0  ��  �:
                �     �Z���� � �����  �  �             ���a�=2    h� �       x  n�  �V
                �     �Z���� � �����  �  �             ���x�W2    o� �       �  0�   s
                �    �Z���� � �����  �  �             ����q2    v� �         �   �
                �    �Z���� � �����  �  �             ��)��2     }� �       P  ��  @�
                �    �Z���� � �����  �  �             ��?��2    (�� �       �  v�  `�
                 �    �Z���� � �����  �  �             ��U�6�2    0�� �       �  8�  ��
   ��            �    �Z���� � �����  �  �             ��k�O�2    8��       (  ��  ��
   ��            �    �Z���� � �����  �  �             ���h�2    @��       p  ��  �   ��   	         �    �Z����    �  �  �              ��i��  2    � � J >         �-  �                �     E������ � �����  �  �              ��w�� ,2    � � N B       /  |.  \�               �     E������ � �����  �  �              ����	82    � � R F       D  l/  ̪               �     E������ � �����  �  �              ����D2    � V J       Z  \0  <�               �    E������ � �����  �  �              ����P2    	� Z N       o  L1  ��               �    E������ � �����  �  �              ����*\2    � ^ R       �  <2  �               �    E������ � �����  �  �              ����5h2    � b V       �  ,3  ��               �    E������ � �����  �  �              ����@t2    � f Z       �  4  ��               �    E������ � �����  �  �              ���K�2    !� j ^       �  5  l�               �    E������ � �����  �  �              ���V�2    '� n b       �  �5  ��   
    	        �    E������ � �����  �  �             ����3m2    � Y M       �  �9  XA                 �     �������	 � �����  �  �             ���?z2    � ] Q       �  �:  �K                �     �������	 � �����  �  �             ���K�2    � a U       �  �;  pV                �     �������	 � �����  �  �             ���*W�2    %� e Y         �<  �`                �    �������	 � �����  �  �             ��;c�2    ,� i ]       2  �=  �k                �    �������	 � �����  �  �             ��Lo�2    3� m a       M  ?  v                �    �������	 � �����  �  �             ��']{�2    :� q e       h  @  ��                �    �������	 � �����  �  �             ��7n��2    A� u i       �  A  ,�                �    �������	 � �����  �  �             ��G��2    H� y m       �  ,B  ��   	             �    �������	 � �����  �  �             ��W���2    O� } q       �  :C  D�        	        �    �������	 � �����  �  �             ��4qx�2    8� h \       �  rG  �      !          �     ۮ�����
 � �����  �  �             ��F���2    ?� l `       �  �H  �      !         �     ۮ�����
 � �����  �  �             ��X���2    F� p d         �I  �+      !         �     ۮ�����
 � �����  �  �             ��j���2    M� t h       >  �J  �8      !         �    ۮ�����
 � �����  �  �             ��|���2    T� x l       _  "L  vE      !         �    ۮ�����
 � �����  �  �             �����2    [� | p       �  NM  ZR      !         �    ۮ�����
 � �����  �  �             �����2    b� � t       �  zN  >_   
   !         �    ۮ�����
 � �����  �  �             �����!2    i� � x       �  �O  "l   	   !         �    ۮ�����
 � �����  �  �             ����/2    p� � |       �  �P  y      !         �    ۮ�����
 � �����  �  �             ����=2    w� �       	  �Q  �      ! 	        �    ۮ�����
 � �����  �  �             �����2    _� v j       f
  �V  (      "           �     E������ � �����  �  �             ����%2    f� { o       �
  �W  �      "          �     E������ � �����  �  �             ����52    m� � t       �
  BY  /      "          �     E������ � �����  �  �             ���+�E2    t� � y       �
  �Z  �>      "          �    E������ � �����  �  �             ���?U2    {� ~         �[  N      "          �    E������ � �����  �  �             ��Se2    �	� �       ,   ]  �]   	   "          �    E������ � �����  �  �             ��!g%u2    �� �       T  j^  �l      "          �    E������ � �����  �  �             ��4{4�2    �� �       |  �_  p|      "          �    E������ � �����  �  �             ��G�C�2    �� �       �  �`  �      "          �    E������ � �����  �  �             ��Z�R�2    �!� �       �  Hb  `�      " 	         �    E������ � �����  �  �             ��.|"z2    �	� �       r  pg  �@      #       !   �     �}Y���� � �����  �  �             ��C�2�2    �� �       �  �h  �R      #      !   �     �}Y���� � �����  �  �             ��X�B�2    �� �       �  @j  @e      #      !   �     �}Y���� � �����  �  �             ��m�R�2    �� �       �  �k  �w   
   #      !   �    �}Y���� � �����  �  �             ����b�2    �!� �       -  m  Љ   	   #      !   �    �}Y���� � �����  �  �             ����r�2    �'� �       \  xn  �      #      !   �    �}Y���� � �����  �  �             ��� ��2    �-� �       �  �o  `�      #      !   �    �}Y���� � �����  �  �             �����2    �3� �       �  Hq  ��      #      !   �    �}Y���� � �����  �  �             ���,�2    �9� �       �  �r  ��      #      !   �    �}Y���� � �����  �  �             ���B�2    �?� �         t  8�      # 	     !   �    �}Y���� � 3   �  �  �             ���}�2    �&� �       
  �y  �      $       "   �     P�b���� � �����  �  �             ���/��2    �,� �       A  >{  d�      $      "   �     P�b���� � �����  �  �             ���G�	2    �2� �       w  �|  ��   	   $      "   �     P�b���� � �����  �  �             �� _�2    �8� �       �  J~  �      $      "   �    P�b���� � �����  �  �             ��w�/2    �>� �       �  �  `�      $      "   �    P�b���� � �����  �  �             ��.��B2    �D� �         V�  �      $      "   �    P�b���� � �����  �  �             ��E��U2    �J� �       R  ܂  (      $      "   �    P�b���� � �����  �  �             ��\��h2    �P� �       �  b�  \=      $      "   �    P�b���� � �����  �  �             ��s�{2    �V� �       �  �  �R      $      "   �    P�b���� � �����  �  �             �����2    �\� �       �  n�  h       $ 	     "   �    P�b���� � 3   �  �  �             ��W��[2    �C� �       :  ��  �J   
   %       #   �     66����� � �����  �  �             ��o��o2    �J� �       y  *�  vc   	   %      #   �     66����� � �����  �  �             �����2    �Q� �       �  ΐ  |      %      #   �     66����� � �����  �  �             ��� �2    �X� �       �  r�  ��      %      #   �    66����� � �����  �  �             ���%3�2    �_� �       6  �  J�      %      #   �    66����� � �����  �  �             ���>F�2    f� �       u  ��  ��      %      #   �    66����� � �����  �  �             ���WY�2    	m� �       �  ^�  ��      %      #   �    66����� � �����  �  �             ���pl�2    t� �       �  �  �      %      #   �    66����� � �����  �  �             ����2    {� �       2  ��  �	   ��  %      #   �    66����� � �����  �  �             ��/��2    !�� �       q  J�  V(	   ��  % 	     #   �    66����� � =   �  �  �             ���oU�2    i� �         ڢ  �-
      &       $   �     ������ � �����  �  �             ���i�2    p� �       V  ��  �I
      &      $   �     ������ � �����  �  �             ��+�}2    w� �       �  ^�  �e
      &      $   �     ������ � �����  �  �             ��E��2    ~� �       �   �   �
      &      $   �    ������ � �����  �  �             ��_��+2    '�� �       .  �   �
      &      $   �    ������ � �����  �  �             ��y��@2    /�� �       v  ��  @�
      &      $   �    ������ � �����  �  �             ����U2    7�� �       �  f�  `�
       &      $   �    ������ � �����  �  �             ���,�j2    ?�� �         (�  ��
   ��  &      $   �    ������ � �����  �  �             ���G�2    G��       N  �  �   ��  &      $   �    ������ � �����  �  �             ���b	�2    O��       �  ��  �*   ��  & 	     $   �    ������ =   �  �  �              ��)`)`2    � R � F       	  �,  ��      3       1   �     ������� � �����  �  �              ��6m6m2    � V � J         �-  �      3      1   �     ������� � �����  �  �              ��CzCz2    � Z � N       4  �.  x�      3      1   �     ������� � �����  �  �              ��P�P�2    � ^ � R       J  �/  �      3      1   �    ������� � �����  �  �              ��]�]�2    � b � V       _  �0  X�      3      1   �    ������� � �����  �  �              ��j�j�2    � f � Z       u  �1  Ƚ      3      1   �    ������� � �����  �  �              ��w�w�2    � j � ^       �  x2  8�      3      1   �    ������� � �����  �  �              ������2    � n � b       �  h3  ��      3      1   �    ������� � �����  �  �              ������2    � r � f       �  X4  �      3      1   �    ������� � �����  �  �              ������2    � v � j       �  H5  ��   
   3 	     1   �    ������� � �����  �  �             ��}�}�2    � a � U       �  9  P:      4       2   �     u������	 � �����  �  �             ������2    � e � Y       �  :  �D      4      2   �     u������	 � �����  �  �             ������2    � i � ]       �  $;  hO      4      2   �     u������	 � �����  �  �             ������2    � m � a         2<  �Y      4      2   �    u������	 � �����  �  �             ������2    � q � e          @=  �d      4      2   �    u������	 � �����  �  �             ����2    u i       ;  N>  o      4      2   �    u������	 � �����  �  �             ����2    y m       V  \?  �y      4      2   �    u������	 � �����  �  �             ��� � 2    } q       q  j@  $�      4      2   �    u������	 � �����  �  �             ���/�/2    � u       �  xA  ��   	   4      2   �    u������	 � �����  �  �             ���>�>2    � y       �  �B  <�      4 	     2   �    u������	 � �����  �  �             ����2    p d       �  �F  *
      5       3   �     vܒ����
 � �����  �  �             ���-�-2    t h       �  �G        5      3   �     vܒ����
 � �����  �  �             ���=�=2    x l       
  I  �#      5      3   �     vܒ����
 � �����  �  �             ��MM2    | p       +  BJ  �0      5      3   �    vܒ����
 � �����  �  �             ��]]2    � t       L  nK  �=      5      3   �    vܒ����
 � �����  �  �             ��&m&m2     �  x       m  �L  �J      5      3   �    vܒ����
 � �����  �  �             ��6}6}2    &� &|       �  �M  �W   
   5      3   �    vܒ����
 � �����  �  �             ��F�F�2    ,� ,�       �  �N  fd   	   5      3   �    vܒ����
 � �����  �  �             ��V�V�2    2� 2�       �  P  Jq      5      3   �    vܒ����
 � �����  �  �             ��f�f�2    8� 8�       �  JQ  .~      5 	     3   �    vܒ����
 � �����  �  �             ��=�=�2     ~  r       Q
  �U  �      6       4   �     �J����� � �����  �  �             ��N�N�2    '� 'w       x
  DW  0      6      4   �     �J����� � �����  �  �             ��_�_�2    .� .|       �
  �X  �&      6      4   �     �J����� � �����  �  �             ��p�p�2    5� 5�       �
  �Y   6      6      4   �    �J����� � �����  �  �             ������2    <� <�       �
  "[  �E      6      4   �    �J����� � �����  �  �             ������2    C� C�         l\  U   	   6      4   �    �J����� � �����  �  �             ������2    J� J�       >  �]  �d      6      4   �    �J����� � �����  �  �             ����2    Q� Q�       f   _   t      6      4   �    �J����� � �����  �  �             ����2    X� X�       �  J`  x�      6      4   �    �J����� � �����  �  �             ���)�)2    _� _�       �  �a  �      6 	     4   �    �J����� � �����  �  �             ��� � 2    G� G�       [  �f  �7      7       5   �     �V#���� � �����  �  �             ����2    N� N�       �  $h  �I      7      5   �     �V#���� � �����  �  �             ���(�(2    U� U�       �  �i  \      7      5   �     �V#���� � �����  �  �             ���<�<2    \� \�       �  �j  dn   
   7      5   �    �V#���� � �����  �  �             ���P�P2    c� c�         \l  ��   	   7      5   �    �V#���� � �����  �  �             ��dd2    j� j�       E  �m  ��      7      5   �    �V#���� � �����  �  �             ��xx2    q� q�       s  ,o  <�      7      5   �    �V#���� � �����  �  �             ��-�-�2    x� x�       �  �p  ��      7      5   �    �V#���� � �����  �  �             ��@�@�2    � �       �  �q  ��      7      5   �    �V#���� � �����  �  �             ��S�S�2    �� ��          ds  �      7 	     5   �    �V#���� � e   �  �  �             ��!�!�2    m� m�       �  y  8�      8       6   �     ��H���� � �����  �  �             ��5�5�2    t� t�       '  �z  ��      8      6   �     ��H���� � �����  �  �             ��I�I�2    {� {�       ^  |  ��   	   8      6   �     ��H���� � �����  �  �             ��]�]�2    �� ��       �  �}  4�      8      6   �    ��H���� � �����  �  �             ��q�q�2    �� ��       �    ��      8      6   �    ��H���� � �����  �  �             ������2    �� ��         ��  �      8      6   �    ��H���� � �����  �  �             ����2    �� ��       8  (�  0      8      6   �    ��H���� � �����  �  �             ����2    �� ��       o  ��  �3      8      6   �    ��H���� � �����  �  �             ���/�/2    �� ��       �  4�  �H      8      6   �    ��H���� � �����  �  �             ���D�D2    �� ��       �  ��  ,^       8 	     6   �    ��H���� � e   �  �  �             ����2    �� ��         Ҍ  N@   
   9       7   �     <|����� � �����  �  �             ���*�*2    �� ��       ^  v�  �X   	   9      7   �     <|����� � �����  �  �             ���A�A2    �� ��       �  �  �q      9      7   �     <|����� � �����  �  �             ���X�X2    �� ��       �  ��  "�      9      7   �    <|����� � �����  �  �             ���o�o2    �� ��         b�  ��      9      7   �    <|����� � �����  �  �             ����2    �� ��       Z  �  Z�      9      7   �    <|����� � �����  �  �             ��#�#�2    �� ��       �  ��  ��      9      7   �    <|����� � �����  �  �             ��9�9�2    �� ��       �  N�  ��      9      7   �    <|����� � �����  �  �             ��O�O�2    �� ��         �  .	   ��  9      7   �    <|����� � �����  �  �             ��e�e�2    �� ��       V  ��  �	   ��  9 	     7   �    <|����� � o   �  �  �             ��+�+�2    �� ��       �  &�  `"
      :       8   �     ׂ����� � �����  �  �             ��B�B�2    �� ��       9  �  �>
      :      8   �     ׂ����� � �����  �  �             ��Y�Y�2    �� ��       �  ��  �Z
      :      8   �     ׂ����� � �����  �  �             ��p�p�2    �� ��       �  l�  �v
      :      8   �    ׂ����� � �����  �  �             ����2    �� ��         .�  ��
      :      8   �    ׂ����� � �����  �  �             ���%�%2    �� ��       Y  �   �
      :      8   �    ׂ����� � �����  �  �             ���=�=2    �� ��       �  ��   �
       :      8   �    ׂ����� � �����  �  �             ���U�U2    ���       �  t�  @�
   ��  :      8   �    ׂ����� � �����  �  �             ���m�m2    �
��       1  6�  `   ��  :      8   �    ׂ����� � �����  �  �             ������2            y  ��  �   ��  : 	     8   �    ׂ����� o   �  �  �              ��Iv@2    � � J >         P-  З      I       F   �     �gQ���� � �����  �  �              ��V�L2    � � N B       )  @.  @�      I      F   �     �gQ���� � �����  �  �              ��c�+X2    � � R F       ?  0/  ��      I      F   �     �gQ���� � �����  �  �              ��p�7d2    � � V J       T   0   �      I      F   �    �gQ���� � �����  �  �              ��}�Cp2    � Z N       j  1  ��      I      F   �    �gQ���� � �����  �  �              ����O|2    
� ^ R       �   2   �      I      F   �    �gQ���� � �����  �  �              ����[�2    � b V       �  �2  p�      I      F   �    �gQ���� � �����  �  �              ����g�2    � f Z       �  �3  ��      I      F   �    �gQ���� � �����  �  �              ����s�2    � j ^       �  �4  P�      I      F   �    �gQ���� � �����  �  �              �����2    "� n b       �  �5  ��   
   I 	     F   �    �gQ���� � �����  �  �             ����]�2    � Y M       �  �9   ?      J       G   �     n�M����	 � �����  �  �             ����j�2    � ] Q       �  �:  �I      J      G   �     n�M����	 � �����  �  �             ����w�2    � a U       �  �;  T      J      G   �     n�M����	 � �����  �  �             �����2     � e Y         �<  �^      J      G   �    n�M����	 � �����  �  �             �����2    '� i ]       ,  �=  0i      J      G   �    n�M����	 � �����  �  �             ���'��2    .� m a       G  �>  �s      J      G   �    n�M����	 � �����  �  �             ���7��2    5� q e       b  �?  H~      J      G   �    n�M����	 � �����  �  �             ��G��2    <� u i       }  �@  Ԉ      J      G   �    n�M����	 � �����  �  �             ��W��2    C� y m       �  �A  `�   	   J      G   �    n�M����	 � �����  �  �             ��$g�2    J� } q       �  �B  �      J 	     G   �    n�M����	 � �����  �  �             �� G��2    3� h \       �  6G  R      K       H   �     ��j����
 � �����  �  �             ��X��2    :� l `       �  bH  6      K      H   �     ��j����
 � �����  �  �             ��"i�2    A� p d         �I  )      K      H   �     ��j����
 � �����  �  �             ��3z�2    H� t h       8  �J  �5      K      H   �    ��j����
 � �����  �  �             ��D��%2    O� x l       Y  �K  �B      K      H   �    ��j����
 � �����  �  �             ��U��42    V� | p       z  M  �O      K      H   �    ��j����
 � �����  �  �             ��f�C2    ]� � t       �  >N  �\   
   K      H   �    ��j����
 � �����  �  �             ��w�R2    d� � x       �  jO  �i   	   K      H   �    ��j����
 � �����  �  �             ����$a2    k� � |       �  �P  rv      K      H   �    ��j����
 � �����  �  �             ����3p2    r� � �       �  �Q  V�      K 	     H   �    ��j����
 � �����  �  �             ��q�	I2    Z� v j       _
  rV  X      L       I   �     J����� � �����  �  �             ����Z2    a� { o       �
  �W  �      L      I   �     J����� � �����  �  �             ����)k2    h� � t       �
  Y  H,      L      I   �     J����� � �����  �  �             ����9|2    o� � y       �
  PZ  �;      L      I   �    J����� � �����  �  �             ���I�2    v� � ~       �
  �[  8K      L      I   �    J����� � �����  �  �             ���Y�2    }� �       %  �\  �Z   	   L      I   �    J����� � �����  �  �             ���-i�2    �
� �       M  .^  (j      L      I   �    J����� � �����  �  �             ���@y�2    �� �       t  x_  �y      L      I   �    J����� � �����  �  �             ��S��2    �� �       �  �`  �      L      I   �    J����� � �����  �  �             ��f��2    �� �       �  b  ��      L 	     I   �    J����� � �����  �  �             ���>j�2    �� �       j  4g  �=      M       J   �     C����� � �����  �  �             ���S{�2    �
� �       �  �h  �O      M      J   �     C����� � �����  �  �             ��h��2    �� �       �  j  4b      M      J   �     C����� � �����  �  �             ��"}��2    �� �       �  lk  |t   
   M      J   �    C����� � �����  �  �             ��6�� 2    �� �       %  �l  Ć   	   M      J   �    C����� � �����  �  �             ��J��2    �"� �       T  <n  �      M      J   �    C����� � �����  �  �             ��^��$2    �(� �       �  �o  T�      M      J   �    C����� � �����  �  �             ��r��62    �.� �       �  q  ��      M      J   �    C����� � �����  �  �             �����H2    �4� �       �  tr  ��      M      J   �    C����� � �����  �  �             ����Z2    �:� �         �s  ,�      M 	     J   �    C����� � �   �  �  �             ��i��+2    �!� �         |y  Ȥ      N       K   �     �s����� � �����  �  �             ��~��?2    �'� �       8  {  �      N      K   �     �s����� � �����  �  �             �����S2    �-� �       o  �|  p�   	   N      K   �     �s����� � �����  �  �             ���g2    �3� �       �  ~  ��      N      K   �    �s����� � �����  �  �             ���'{2    �9� �       �  �  �      N      K   �    �s����� � �����  �  �             ���=.�2    �?� �         �  l      N      K   �    �s����� � �����  �  �             ���SA�2    �E� �       I  ��  �$      N      K   �    �s����� � �����  �  �             ���iT�2    �K� �       �  &�  :      N      K   �    �s����� � �����  �  �             ��g�2    �Q� �       �  ��  hO      N      K   �    �s����� � �����  �  �             ��&�z�2    �W� �       �  2�  �d       N 	     K   �    �s����� � �   �  �  �             ���eC�2    �>� �       1  J�  VG   
   O       L   �     ��H���� � �����  �  �             ��}W�2    �E� �       p  �  �_   	   O      L   �     ��H���� � �����  �  �             ���k�2    �L� �       �  ��  �x      O      L   �     ��H���� � �����  �  �             ��6��2    �S� �       �  6�  *�      O      L   �    ��H���� � �����  �  �             ��M��2    �Z� �       -  ړ  Ʃ      O      L   �    ��H���� � �����  �  �             ��d��2    �a� �       l  ~�  b�      O      L   �    ��H���� � �����  �  �             ��{��+2    h� �       �  "�  ��      O      L   �    ��H���� � �����  �  �             ����@2    o� �       �  Ƙ  ��      O      L   �    ��H���� � �����  �  �             ���%�U2    v� �       )  j�  6	   ��  O      L   �    ��H���� � �����  �  �             ���=�j2    }� �       h  �  �$	   ��  O 	     L   �    ��H���� � �   �  �  �             ���	�32    d� �         ��  �)
      P       M   �     ������� � �����  �  �             ���#�J2    
k� �       L  `�   F
      P      M   �     ������� � �����  �  �             ���=�a2    r� �       �  "�   b
      P      M   �     ������� � �����  �  �             ���W�x2    y� �       �  �  @~
      P      M   �    ������� � �����  �  �             ���q�2    "�� �       $  ��  `�
      P      M   �    ������� � �����  �  �             ���)�2    *�� �       l  h�  ��
      P      M   �    ������� � �����  �  �             ���?�2    2�� �       �  *�  ��
       P      M   �    ������� � �����  �  �             ��6�U�2    :�� �       �  �  ��
   ��  P      M   �    ������� � �����  �  �             ��O�k�2    B��       D  ��  �
   ��  P      M   �    ������� � �����  �  �             ��h��2    J��       �  p�   '   ��  P 	     M   �    ������� �   �  �  �              ���  i�2    Q  � D       �  `,  `�      _       [   �     ^l����� � �����  �  �              ��� ,w�2    U � � H         P-  З      _      [   �     ^l����� � �����  �  �              ��	8��2    Y � � L       )  @.  @�      _      [   �     ^l����� � �����  �  �              ��D��2    ] � � P       ?  0/  ��      _      [   �    ^l����� � �����  �  �              ��P��2    a � � T       T   0   �      _      [   �    ^l����� � �����  �  �              ��*\��2    e � X       j  1  ��      _      [   �    ^l����� � �����  �  �              ��5h��2    i � \       �   2   �      _      [   �    ^l����� � �����  �  �              ��@t��2    m � `       �  �2  p�      _      [   �    ^l����� � �����  �  �              ��K��2    q � d       �  �3  ��      _      [   �    ^l����� � �����  �  �              ��V��2    u � h       �  �4  P�   
   _ 	     [   �    ^l����� � �����  �  �             ��3m��2    ` � S       �  �8  �5      `       \   �     � ����	 � �����  �  �             ��?z�2    d � W       �  �9  ,@      `      \   �     � ����	 � �����  �  �             ��K��2    h � [       �  �:  �J      `      \   �     � ����	 � �����  �  �             ��W��*2    l � _       �  �;  DU      `      \   �    � ����	 � �����  �  �             ��c�;2    p � "c         �<  �_      `      \   �    � ����	 � �����  �  �             ��o�L2    t � )g       /  �=  \j      `      \   �    � ����	 � �����  �  �             ��{�']2    x � 0k       J  �>  �t      `      \   �    � ����	 � �����  �  �             ����7n2    | � 7o       e  �?  t      `      \   �    � ����	 � �����  �  �             ����G2    � � >s       �   A   �   	   `      \   �    � ����	 � �����  �  �             ����W�2    � � Ew       �  B  ��      ` 	     \   �    � ����	 � �����  �  �             ��x�4q2    o � .b       �  FF        a       ]   �     �\����
 � �����  �  �             ����F�2    t � 5f       �  rG  �      a      ]   �     �\����
 � �����  �  �             ����X�2    y � <j       �  �H  �      a      ]   �     �\����
 � �����  �  �             ����j�2    ~ � Cn         �I  �+      a      ]   �    �\����
 � �����  �  �             ����|�2    � � Jr       >  �J  �8      a      ]   �    �\����
 � �����  �  �             �����2    � � Qv       _  "L  vE      a      ]   �    �\����
 � �����  �  �             �����2    � � Xz       �  NM  ZR   
   a      ]   �    �\����
 � �����  �  �             ���!��2    � � _~       �  zN  >_   	   a      ]   �    �\����
 � �����  �  �             ���/�2    � � f�       �  �O  "l      a      ]   �    �\����
 � �����  �  �             ���=�2    � � m�       �  �P  y      a 	     ]   �    �\����
 � �����  �  �             �����2    � � Up       B
  �U        b       ^   �      l����� � �����  �  �             ���%�2    � � \u       j
  �V  �      b      ^   �      l����� � �����  �  �             ���5�2    � � cz       �
  X  !      b      ^   �      l����� � �����  �  �             ���E�+2    � � j       �
  `Y  �0      b      ^   �     l����� � �����  �  �             ��U�?2    � � q�       �
  �Z  �?      b      ^   �     l����� � �����  �  �             ��eS2    � � x�         �[  pO   	   b      ^   �     l����� � �����  �  �             ��%u!g2    � � �       0  >]  �^      b      ^   �     l����� � �����  �  �             ��4�4{2    � � ��       X  �^  `n      b      ^   �     l����� � �����  �  �             ��C�G�2    � � ��         �_  �}      b      ^   �     l����� � �����  �  �             ��R�Z�2    � � ��       �  a  P�      b 	     ^   �     l����� � �����  �  �             ��"z.|2    � � {�       K  Df  t1      c       _   �     Cc���� � �����  �  �             ��2�C�2    � � ��       z  �g  �C      c      _   �     Cc���� � �����  �  �             ��B�X�2    � � ��       �  i  V      c      _   �     Cc���� � �����  �  �             ��R�m�2    � � ��       �  |j  Lh   
   c      _   �    Cc���� � �����  �  �             ��b���2    � � ��         �k  �z   	   c      _   �    Cc���� � �����  �  �             ��r���2    �  ��       5  Lm  ܌      c      _   �    Cc���� � �����  �  �             ����� 2    � ��       d  �n  $�      c      _   �    Cc���� � �����  �  �             �����2    � ��       �  p  l�      c      _   �    Cc���� � �����  �  �             ����,2    � ��       �  �q  ��      c      _   �    Cc���� � �����  �  �             ����B2    � ��       �  �r  ��      c 	     _   �    Cc���� � �   �  �  �             ��}��2    �  ��       �  �x  ��      d       `   �     Y#V���� � �����  �  �             �����/2    � ��         z  ��      d      `   �     Y#V���� � �����  �  �             ���	�G2    � ��       M  �{  P�   	   d      `   �     Y#V���� � �����  �  �             ��� _2    � ��       �  }  ��      d      `   �    Y#V���� � �����  �  �             ���/w2    � ��       �  �~  ��      d      `   �    Y#V���� � �����  �  �             ���B.�2    � ��       �  *�  L      d      `   �    Y#V���� � �����  �  �             ���UE�2    � $��       (  ��  �      d      `   �    Y#V���� � �����  �  �             ���h\�2    � *��       ^  6�  �,      d      `   �    Y#V���� � �����  �  �             ��{s�2    � 0��       �  ��  HB      d      `   �    Y#V���� � �����  �  �             �����2    � 6��       �  B�  �W       d 	     `   �    Y#V���� � �   �  �  �             ���[W�2    � ��         Z�  F9   
   e       a   �     �y ���� � �����  �  �             ���oo�2    � $��       L  ��  �Q   	   e      a   �     �y ���� � �����  �  �             �����2    � *��       �  ��  ~j      e      a   �     �y ���� � �����  �  �             �� ��2    � 0��       �  F�  �      e      a   �    �y ���� � �����  �  �             ��3��%2    � 6��       	  �  ��      e      a   �    �y ���� � �����  �  �             ��F��>2    � <��       H  ��  R�      e      a   �    �y ���� � �����  �  �             ��Y��W2    � B��       �  2�  ��      e      a   �    �y ���� � �����  �  �             ��l��p2    � H�       �  ֗  ��      e      a   �    �y ���� � �����  �  �             ����2    � N�         z�  &�   ��  e      a   �    �y ���� � �����  �  �             ���/�2    T�       D  �  �	   ��  e 	     a   �    �y ���� � �   �  �  �             ��U��o2    � ;��       �  ��  �
      f       b   �     ������ � �����  �  �             ��i��2    � B�       &  p�   7
      f      b   �     ������ � �����  �  �             ��}+�2    � I�       n  2�   S
      f      b   �     ������ � �����  �  �             ���E�2    � P�       �  ��  @o
      f      b   �    ������ � �����  �  �             ���+_�2    W�       �  ��  `�
      f      b   �    ������ � �����  �  �             ���@y�2    ^%�       F  x�  ��
      f      b   �    ������ � �����  �  �             ���U�2    e-�       �  :�  ��
       f      b   �    ������ � �����  �  �             ���j�,2    l5�       �  ��  ��
   ��  f      b   �    ������ � �����  �  �             ����G2    s=�         ��  ��
   ��  f      b   �    ������ � �����  �  �             ��	��b2    #zE      f  ��      ��  f 	     b   �    ������ �   �  �  �               KK
2    � R � F         -  ��      y       s   �     ������� � �����  �  �               *X*X
2    � V � J       $  .  $�      y      s   �     ������� � �����  �  �               6e6e
2    � Z � N       9  �.  ��      y      s   �     ������� � �����  �  �               BrBr
2    � ^ � R       O  �/  �      y      s   �    ������� � �����  �  �               NN
2    � b � V       e  �0  t�      y      s   �    ������� � �����  �  �               Z�Z�
2    � f � Z       z  �1  �      y      s   �    ������� � �����  �  �               f�f�
2    � j � ^       �  �2  T�      y      s   �    ������� � �����  �  �               r�r�
2    � n � b       �  �3  ��      y      s   �    ������� � �����  �  �               ~�~�
2    � r � f       �  �4  4�      y      s   �    ������� � �����  �  �               ����
2    � v � j       �  �5  ��   
   y 	     s   �    ������� � �����  �  �              h�h�
2    � a � U       �  D9  �<      z       t   �     �������	 � �����  �  �              v�v�
2    � e � Y       �  R:  4G      z      t   �     �������	 � �����  �  �              ����
2    � i � ]       �  `;  �Q      z      t   �     �������	 � �����  �  �              ����
2    � m � a         n<  L\      z      t   �    �������	 � �����  �  �              ����
2    � q � e       &  |=  �f      z      t   �    �������	 � �����  �  �              ����
2    � u i       A  �>  dq      z      t   �    �������	 � �����  �  �              ����
2    y m       \  �?  �{      z      t   �    �������	 � �����  �  �              ��
2    } q       w  �@  |�      z      t   �    �������	 � �����  �  �              ��
2    � u       �  �A  �   	   z      t   �    �������	 � �����  �  �              � � 
2    � y       �  �B  ��      z 	     t   �    �������	 � �����  �  �              ����
2     p d       �  �F  �      {       u   �     �������
 � �����  �  �              ��
2    t h       �  &H  �      {      u   �     �������
 � �����  �  �              ��
2    x l         RI  �&      {      u   �     �������
 � �����  �  �              �.�.
2    | p       1  ~J  j3      {      u   �    �������
 � �����  �  �              �>�>
2    � t       R  �K  N@      {      u   �    �������
 � �����  �  �              NN
2    �  x       s  �L  2M      {      u   �    �������
 � �����  �  �              ^^
2    $� &|       �  N  Z   
   {      u   �    �������
 � �����  �  �              *n*n
2    *� ,�       �  .O  �f   	   {      u   �    �������
 � �����  �  �              9~9~
2    0� 2�       �  ZP  �s      {      u   �    �������
 � �����  �  �              H�H�
2    6� 8�       �  �Q        { 	     u   �    �������
 � �����  �  �              hh
2    ~  r       X
  6V  �
      |       v   �     ������� � �����  �  �              /y/y
2    %� 'w       �
  �W         |      v   �     ������� � �����  �  �              @�@�
2    ,� .|       �
  �X  x)      |      v   �     ������� � �����  �  �              Q�Q�
2    3� 5�       �
  Z  �8      |      v   �    ������� � �����  �  �              b�b�
2    :� <�       �
  ^[  hH      |      v   �    ������� � �����  �  �              s�s�
2    A� C�         �\  �W   	   |      v   �    ������� � �����  �  �              ����
2    H� J�       F  �]  Xg      |      v   �    ������� � �����  �  �              ����
2    O� Q�       m  <_  �v      |      v   �    ������� � �����  �  �              ����
2    V� X�       �  �`  H�      |      v   �    ������� � �����  �  �              ��
2    ]� _�       �  �a  ��      | 	     v   �    ������� � �����  �  �              ����
2    E� G�       b  �f  �:      }       w   �     ������� � �����  �  �              ����
2    L� N�       �  `h  �L      }      w   �     ������� � �����  �  �              ����
2    S� U�       �  �i  (_      }      w   �     ������� � �����  �  �              ��
2    Z� \�       �  0k  pq   
   }      w   �    ������� � �����  �  �              �#�#
2    a� c�         �l  ��   	   }      w   �    ������� � �����  �  �              �6�6
2    h� j�       L   n   �      }      w   �    ������� � �����  �  �              �I�I
2    o� q�       {  ho  H�      }      w   �    ������� � �����  �  �              \\
2    v� x�       �  �p  ��      }      w   �    ������� � �����  �  �              oo
2    }� �       �  8r  ��      }      w   �    ������� � �����  �  �              +�+�
2    �� ��         �s   �      } 	     w   �    ������� � �   �  �  �              �T�T
2    k� m�       �  @y  ��      ~       x   �     ������� � �����  �  �              hh
2    r� t�       0  �z  Զ      ~      x   �     ������� � �����  �  �              ||
2    y� {�       f  L|  (�   	   ~      x   �     ������� � �����  �  �              1�1�
2    �� ��       �  �}  |�      ~      x   �    ������� � �����  �  �              D�D�
2    �� ��       �  X  ��      ~      x   �    ������� � �����  �  �              W�W�
2    �� ��       
  ހ  $      ~      x   �    ������� � �����  �  �              j�j�
2    �� ��       A  d�  x!      ~      x   �    ������� � �����  �  �              }�}�
2    �� ��       w  �  �6      ~      x   �    ������� � �����  �  �              ����
2    �� ��       �  p�   L      ~      x   �    ������� � �����  �  �              ��
2    �� ��       �  ��  ta       ~ 	     x   �    ������� � �   �  �  �              l�l�
2    �� ��       (  �  �C   
          y   �     ������� � �����  �  �              ����
2    �� ��       g  ��  n\   	         y   �     ������� � �����  �  �              ��
2    �� ��       �  V�  
u            y   �     ������� � �����  �  �              ��
2    �� ��       �  ��  ��            y   �    ������� � �����  �  �              �.�.
2    �� ��       $  ��  B�            y   �    ������� � �����  �  �              �D�D
2    �� ��       c  B�  ޾            y   �    ������� � �����  �  �              �Z�Z
2    �� ��       �  �  z�            y   �    ������� � �����  �  �              �p�p
2    �� ��       �  ��  �            y   �    ������� � �����  �  �              ��
2    �� ��          .�  �	   ��        y   �    ������� � �����  �  �              )�)�
2    �� ��       _  қ  N!	   ��   	     y   �    ������� �   �  �  �              �f�f
2    �� ��       �  b�   &
      �       z   �     ������� � �����  �  �              }}
2    �� ��       C  $�  @B
      �      z   �     ������� � �����  �  �              ��
2    �� ��       �  �  `^
      �      z   �     ������� � �����  �  �              0�0�
2    �� ��       �  ��  �z
      �      z   �    ������� � �����  �  �              F�F�
2    �� ��         j�  ��
      �      z   �    ������� � �����  �  �              \�\�
2    �� ��       c  ,�  ��
      �      z   �    ������� � �����  �  �              r�r�
2    �� ��       �  �  ��
       �      z   �    ������� � �����  �  �              ��
2    ���       �  ��   �
   ��  �      z   �    ������� � �����  �  �              ��
2    �
��       ;  r�      ��  �      z   �    ������� � �����  �  �              �5�5
2    �       �  4�  @#   ��  � 	     z   �    �������   �  �  �              ��\��  2    � � J >         �-  �       �       �   �     ���������� �����  �  �              ��j�� ,2    � � N B       4  �.  x�       �      �   �     ���������� �����  �  �              ��x�	82    � � R F       J  �/  �       �      �   �     ���������� �����  �  �              ����D2    � � V J       _  �0  X�       �      �   �    ���������� �����  �  �              ����P2    � � Z N       u  �1  Ƚ       �      �   �    ���������� �����  �  �              ����*\2    � � ^ R       �  x2  8�       �      �   �    ���������� �����  �  �              ����5h2    � � b V       �  h3  ��       �      �   �    ���������� �����  �  �              ����@t2    � � f Z       �  X4  �       �      �   �    ���������� �����  �  �              ���K�2    � � j ^       �  H5  ��       �      �   �    ���������� �����  �  �              ���V�2    � n b       �  86  ��       � 	     �   �    ���������� �����  �  �             ����3m2    � � Y M       �  �9  �C       �       �   �     ���������� �����  �  �             ���?z2    � � ] Q       �  ;  <N       �      �   �     ���������� �����  �  �             ���K�2    � � a U         <  �X       �      �   �     ���������� �����  �  �             ���$W�2    � � e Y         "=  Tc       �      �   �    ���������� �����  �  �             ���4c�2    � i ]       8  0>  �m       �      �   �    ���������� �����  �  �             ��Do�2    	m a       S  >?  lx       �      �   �    ���������� �����  �  �             ��T{�2    
q e       n  L@  ��       �      �   �    ���������� �����  �  �             ��#d��2    u i       �  ZA  ��       �      �   �    ���������� �����  �  �             ��2t��2    y m       �  hB  �       �      �   �    ���������� �����  �  �             ��A���2    !} q       �  vC  ��       � 	     �   �    ���������� �����  �  �             ��dx�2    
h \       �  �G  z       �       �   �     ���������� �����  �  �             ��.v��2    l `         �H  ^!       �      �   �     ���������� �����  �  �             ��?���2    p d       $  J  B.       �      �   �     ���������� �����  �  �             ��P���2    t h       E  2K  &;       �      �   �    ���������� �����  �  �             ��a���2    "x l       f  ^L  
H       �      �   �    ���������� �����  �  �             ��r��2    (#| p       �  �M  �T       �      �   �    ���������� �����  �  �             �����2    .)� t       �  �N  �a       �      �   �    ���������� �����  �  �             �����!2    4/� x       �  �O  �n       �      �   �    ���������� �����  �  �             �����/2    :5� |       �  Q  �{       �      �   �    ���������� �����  �  �             ����=2    @;� �       	  :R  ~�       � 	     �   �    ���������� �����  �  �             �����2    (#v j       n
  �V  �       �       �        ���������� �����  �  �             �����%2    /*{ o       �
  4X  p"       �      �        ���������� �����  �  �             ���
�52    61� t       �
  ~Y  �1       �      �        ���������� �����  �  �             ����E2    =8� y       �
  �Z  `A       �      �       ���������� �����  �  �             ���2U2    D?� ~         \  �P       �      �       ���������� �����  �  �             ���Fe2    KF� �       4  \]  P`       �      �       ���������� �����  �  �             �� Z%u2    RM� �       [  �^  �o       �      �       ���������� �����  �  �             ��n4�2    YT� �       �  �_  @       �      �       ���������� �����  �  �             ��&�C�2    `[� �       �  :a  ��       �      �       ���������� �����  �  �             ��9�R�2    gb� �       �  �b  0�       � 	     �       ���������� �����  �  �             ��o"z2    OJ� �       z  �g  �C       �       �       ���������� �����  �  �             ��!�2�2    VQ� �       �  i  V       �      �       ���������� �����  �  �             ��5�B�2    ]X� �       �  |j  Lh       �      �       ���������� �����  �  �             ��I�R�2    d_� �         �k  �z       �      �      ���������� �����  �  �             ��]�b�2    kf� �       5  Lm  ܌       �      �      ���������� �����  �  �             ��q�r�2    rm� �       d  �n  $�       �      �      ���������� �����  �  �             ������2    yt� �       �  p  l�       �      �      ���������� �����  �  �             �����2    �{� �       �  �q  ��       �      �      ���������� �����  �  �             ����2    ��� �       �  �r  ��       �      �      ���������� �����  �  �             ���,�2    ��� �         Tt  D�       � 	     �      ���������� �����  �  �             ��� }�2    up� �         �y  X�       �       �       ���������� �����  �  �             �����2    |w� �       I  z{  ��       �      �       ���������� �����  �  �             ���.�	2    �~� �       �   }   �       �      �       ���������� �����  �  �             ���E�2    ��� �       �  �~  T�       �      �      ���������� �����  �  �             ���\�/2    ��� �       �  �  �        �      �      ���������� �����  �  �             ���s�B2    ��� �       #  ��  �       �      �      ���������� �����  �  �             ����U2    ��� �       Z  �  P+       �      �      ���������� �����  �  �             ��*��h2    ��� �       �  ��  �@       �      �      ���������� �����  �  �             ��@�{2    ��� �       �  $�  �U       �      �      ���������� �����  �  �             ��V��2    ��� �       �  ��  Lk       � 	     �      ���������� �����  �  �             ��"��[2    ��� �       C    ^N       �       �       ���������� �����  �  �             ��:��o2    ��� �       �  f�  �f       �      �       ���������� �����  �  �             ��R��2    ��� �       �  
�  �       �      �       ���������� �����  �  �             ��j� �2    ��� �          ��  2�       �      �      ���������� �����  �  �             ���3�2    ��� �       ?  R�  ΰ       �      �      ���������� �����  �  �             ���F�2    ��� �       ~  ��  j�       �      �      ���������� �����  �  �             ���6Y�2    ��� �       �  ��  �       �      �      ���������� �����  �  �             ���Ol�2    ��� �       �  >�  ��       �      �      ���������� �����  �  �             ���h�2    ��� �       ;  �  >	       �      �      ���������� �����  �  �             �����2    ��� �       z  ��  �+	       � 	     �      ���������� �����  �  �             ���NU�2    ��� �         �  `1
       �       �       ���������� �����  �  �             ���ii�2    ��� �       `  ؤ  �M
       �      �       ���������� �����  �  �             ����}2    ��� �       �  ��  �i
       �      �       ���������� �����  �  �             ����2    ��� �       �  \�  ��
       �      �      ���������� �����  �  �             ��&��+2    ��� �       8  �  �
       �      �      ���������� �����  �  �             ��?��@2    ��� �       �  �   �
       �      �      ���������� �����  �  �             ��X��U2    ��� �       �  ��   �
       �      �      ���������� �����  �  �             ��q�j2    ��� �         d�  @�
       �      �      ���������� �����  �  �             ���&�2     ��       X  &�  `       �      �      ���������� �����  �  �             ���A	�2    �       �  �  �.       � 	     �      ��������������  �  �           ����              � T - !         \  (n               ��        ���� � �������������          ����              � X 0 $       #  �  �q              ��        ���� � �������������          ����              � \ 3 '       ,  �  0u              ��        ���� � �������������          ����     !          � ` 6 *       5    �x              ��       ���� � �������������          ����   " #          � d 9 -       >  �  8|              ��       ���� � �������������          ����   $ %          � h < 0       G  J  �              ��       ���� � �������������          ����   & '          � l ? 3       P  �  @�              ��       ���� � �������������          ����   ( )          � p B 6       Y  v  Ć              ��       ���� � �������������          ����   + ,          � t E 9       b    H�    
          ��       ���� � �������������          ����   - .          � x H <       k  �  ̍    	   	       ��       ���� � �������������           ����              � c 4 (       �  �  ֵ               ��        ���� � �������������          ����     !          � h 7 +       �  �  º              ��        ���� � �������������          ����   " #          � m : .       �  b  ��              ��        ���� � �������������          ����   % &          � r = 1       �    ��              ��       ���� � �������������          ����   ' (          � w @ 4         �  ��              ��       ���� � �������������          ����   ) *          � | C 7         ~  r�              ��       ���� � �������������          ����   + ,          � � F :         2  ^�              ��       ���� � �������������          ����   - .          � � I =       )  �  J�    	          ��       ���� � �������������          ����   0 1          � � L @       6  �  6�              ��       ���� � �������������          ����   2 3          � � O C       B  N   "�       	       ��       ���� � �������������          ����   # $          � { : .       �  #  �              ��        ���� � �����  �  �          ����   % &          � � > 2       �  �#  �             ��        ���� � �����  �  �          ����   ' (          � � B 6       �  �$  &             ��        ���� � �����  �  �          ����   * +          � � F :         �%  �,             ��       ���� � �����  �  �          ����   , -          � J >         f&  03             ��       ���� � �����  �  �          ����   . /          � N B       #  8'  �9   	          ��       ���� � �����  �  �          ����   0 1          � R F       4  
(  P@             ��       ���� � �����  �  �          ����   2 3          � V J       D  �(  �F             ��       ���� � �����  �  �          ����   5 6          � Z N       U  �)  pM             ��       ���� � �����  �  �          ����   7 8          � ^ R       f  �*   T      	       ��       ���� � �����  �  �          ����   ( )          	� J >         �-  �              ��        ���� � �����  �  �          ����   * +          � N B       4  �.  x�             ��        ���� � �����  �  �          ����   , -          � R F       J  �/  �             ��        ���� � �����  �  �          ����   / 0          � V J       _  �0  X�   	          ��       ���� � �����  �  �          ����   1 2          %� Z N       u  �1  Ƚ             ��       ���� � �����  �  �          ����   3 4          ,� ^ R       �  x2  8�             ��       ���� � �����  �  �          ����   5 6          3� b V       �  h3  ��             ��       ���� � �����  �  �          ����   7 8          :� f Z       �  X4  �             ��       ���� � �����  �  �          ����   : ;          A� j ^       �  H5  ��             ��       ���� � �����  �  �          ����   < =          H� n b       �  86  ��      	       ��       ���� � -  �  �  �          ����   - .          2� Y M       �  �9  �C            	  ��	        ����	 � �����  �  �          ����   / 0          9� ] Q       �  ;  <N   
        	  ��	        ����	 � �����  �  �          ����   1 2          @� a U         <  �X           	  ��	        ����	 � �����  �  �          ����   4 5          G� e Y         "=  Tc           	  ��	       ����	 � �����  �  �          ����   6 7          N� i ]       8  0>  �m           	  ��	       ����	 � �����  �  �          ����   8 9          U� m a       S  >?  lx           	  ��	       ����	 � �����  �  �          ����   : ;          \� q e       n  L@  ��           	  ��	       ����	 � �����  �  �          ����   < =          c� u i       �  ZA  ��           	  ��	       ����	 � �����  �  �          ����   ? @          j� y m       �  hB  �            	  ��	       ����	 � �����  �  �          ����   A B          q� } q       �  vC  ��   ��  	     	  ��	       ����	 � 7  �  �  �           ����              A ^ � '         \  (n       .        ��
        ���� � �������������          ����              D b � *       #  �  �q       .       ��
        ���� � �������������          ����              G f � -       ,  �  0u       .       ��
        ���� � �������������          ����              J j � 0       5    �x       .       ��
       ���� � �������������          ����              M n � 3       >  �  8|       .       ��
       ���� � �������������          ����              P r � 6       G  J  �       .       ��
       ���� � �������������          ����     !          S v � 9       P  �  @�       .       ��
       ���� � �������������          ����   " #          V z � <       Y  v  Ć       .       ��
       ���� � �������������          ����   $ %          Y ~ � ?       b    H�    
   .       ��
       ���� � �������������          ����   & '          \ � � B       k  �  ̍    	   .	       ��
       ���� � �������������           ����              H m � .       �  �  ֵ       /        ��        ���� � �������������          ����              L q � 1       �  �  º       /       ��        ���� � �������������          ����              P u � 4       �  b  ��       /       ��        ���� � �������������          ����              T y � 7       �    ��       /       ��       ���� � �������������          ����               X } � :         �  ��       /       ��       ���� � �������������          ����   " #          \ � � =         ~  r�       /       ��       ���� � �������������          ����   $ %          ` � � @         2  ^�       /       ��       ���� � �������������          ����   & '          d � � C       )  �  J�    	   /       ��       ���� � �������������          ����   ( )          h � � F       6  �  6�       /       ��       ���� � �������������          ����   * +          l � � I       B  N   "�       /	       ��       ���� � �������������          ����              X | � 4       �  #  �      0        ��        ���� � �����  �  �          ����              \ � � 8       �  �#  �      0       ��        ���� � �����  �  �          ����               ` � � <       �  �$  &      0       ��        ���� � �����  �  �          ����   ! "          d � � @         �%  �,      0       ��       ���� � �����  �  �          ����   # $          h � � D         f&  03      0       ��       ���� � �����  �  �          ����   % &          l �  H       #  8'  �9   	   0       ��       ���� � �����  �  �          ����   ( )          p � L       4  
(  P@      0       ��       ���� � �����  �  �          ����   * +          t � P       D  �(  �F      0       ��       ���� � �����  �  �          ����   , -          x � T       U  �)  pM      0       ��       ���� � �����  �  �          ����   . /          | � X       f  �*   T      0	       ��       ���� � �����  �  �          ����               h � D         �-  �      1        ��        ���� � �����  �  �          ����   ! "          l � 	H       4  �.  x�      1       ��        ���� � �����  �  �          ����   # $          p � L       J  �/  �      1       ��        ���� � �����  �  �          ����   % &          t � P       _  �0  X�   	   1       ��       ���� � �����  �  �          ����   ' (          x � T       u  �1  Ƚ      1       ��       ���� � �����  �  �          ����   ) *          | � %X       �  x2  8�      1       ��       ���� � �����  �  �          ����   , -          � � ,\       �  h3  ��      1       ��       ���� � �����  �  �          ����   . /          � � 3`       �  X4  �      1       ��       ���� � �����  �  �          ����   0 1          � � :d       �  H5  ��      1       ��       ���� � �����  �  �          ����   2 3          � � Ah       �  86  ��      1	       ��       ���� � -  �  �  �          ����   # $          w � +S       �  �9  �C      2      	  ��        ����	 � �����  �  �          ����   % &          { � 2W       �  ;  <N   
   2     	  ��        ����	 � �����  �  �          ����   ' (           � 9[         <  �X      2     	  ��        ����	 � �����  �  �          ����   ) *          � � @_         "=  Tc      2     	  ��       ����	 � �����  �  �          ����   + ,          � � Gc       8  0>  �m      2     	  ��       ����	 � �����  �  �          ����   - .          � � Ng       S  >?  lx      2     	  ��       ����	 � �����  �  �          ����   0 1          � � Uk       n  L@  ��      2     	  ��       ����	 � �����  �  �          ����   2 3          � � \o       �  ZA  ��      2     	  ��       ����	 � �����  �  �          ����   4 5          � � cs       �  hB  �       2     	  ��       ����	 � �����  �  �          ����   6 7          � � jw       �  vC  ��   ��  2	     	  ��       ����	 � 7  �  �  �           ����              .   .         	      �       >        ��        ���� � �������������           ����              2   2            >  |       >       ��        ���� � �������������           ����              6   6            \  �       >       ��        ���� � �������������           ����    	          :   :            z  �       >       ��       ���� � �������������           ����   
           >   >            �  0       >       ��       ���� � �������������           ����              B   B            �  l       >       ��       ���� � �������������           ����              F   F            �  �       >       ��       ���� � �������������           ����              J   J            �  �       >       ��       ���� � �������������           ����              N   N                      >       ��       ���� � �������������           ����              R   R            .  \       >	       ��       ���� � �������������           ����              @  @         #   �  �       ?        ��        ���� � �������������           ����    	          D  D         %   �  �       ?       ��        ���� � �������������           ����   
           H  H         '     Z       ?       ��        ���� � �������������           ����              L  L         )   Z         ?       ��       ���� � �������������           ����              P  P         *   �  �       ?       ��       ���� � �������������           ����              T  T         ,   �  v       ?       ��       ���� � �������������           ����              X  X         .     *       ?       ��       ���� � �������������           ����              \ ! \         0   J  �       ?       ��       ���� � �������������           ����              ` # `         2   �  �       ?       ��       ���� � �������������           ����              d % d         3   �  F       ?	       ��       ���� � �������������           ����   
           Q  Q        N   �  �       @        ��        ���� � �������������          ����              V  V        R     0        @       ��        ���� � �������������          ����              [  [        V   f  �!       @       ��        ���� � �������������          ����              `  `        Y   �   #       @       ��       ���� � �������������          ����              e  e        ]   	  h$       @       ��       ���� � �������������          ����              j   j "       `   t	  �%       @       ��       ���� � �������������          ����              o # o %       d   �	  8'       @       ��       ���� � �������������          ����              t & t (       h   (
  �(       @       ��       ���� � �������������          ����              y ) y +       k   �
  *       @       ��       ���� � �������������          ����              ~ , ~ .       o   �
  p+       @	       ��       ���� � �������������           ����              k  k        �   D  T=       A        ��        ���� � �������������          ����              p  p        �   �  �?       A       ��        ���� � �������������          ����              u  u !       �   4  B       A       ��        ���� � �������������          ����              z " z $       �   �  \D       A       ��       ���� � �������������          ����               %  '       �   $  �F       A       ��       ���� � �������������          ����              � ( � *       �   �  I       A       ��       ���� � �������������          ����              � + � -       �     dK       A       ��       ���� � �������������          ����              � . � 0       �   �  �M       A       ��       ���� � �������������          ����               � 1 � 3       �     P       A       ��       ���� � �������������          ����   ! "          � 4 � 6       �   |  lR       A	       ��       ���� � �������������           ����              �   � "         \  (n       B        ��        ���� � �������������          ����              � # � %       #  �  �q       B       ��        ���� � �������������          ����              � & � (       ,  �  0u       B       ��        ���� � �������������          ����              � ) � +       5    �x       B       ��       ���� � �������������          ����              � , � .       >  �  8|       B       ��       ���� � �������������          ����              � / � 1       G  J  �       B       ��       ���� � �������������          ����               � 2 � 4       P  �  @�       B       ��       ���� � �������������          ����   ! "          � 5 � 7       Y  v  Ć       B       ��       ���� � �������������          ����   # $          � 8 � :       b    H�    
   B       ��       ���� � �������������          ����   % &          � ; � =       k  �  ̍    	   B	       ��       ���� � �������������           ����              � ' � )       �  �  ֵ       C        ��        ���� � �������������          ����              � * � ,       �  �  º       C       ��        ���� � �������������          ����              � - � /       �  b  ��       C       ��        ���� � �������������          ����              � 0 � 2       �    ��       C       ��       ���� � �������������          ����              � 3 � 5         �  ��       C       ��       ���� � �������������          ����   ! "          � 6 � 8         ~  r�       C       ��       ���� � �������������          ����   # $          � 9 � ;         2  ^�       C       ��       ���� � �������������          ����   % &          � < � >       )  �  J�    	   C       ��       ���� � �������������          ����   ' (          � ? � A       6  �  6�       C       ��       ���� � �������������          ����   ) *          � B � D       B  N   "�       C	       ��       ���� � �������������          ����              � - � /       �  #  �      D        ��        ���� � �����  �  �          ����              � 1 � 3       �  �#  �      D       ��        ���� � �����  �  �          ����              � 5 � 7       �  �$  &      D       ��        ���� � �����  �  �          ����     !          � 9 � ;         �%  �,      D       ��       ���� � �����  �  �          ����   " #          � = � ?         f&  03      D       ��       ���� � �����  �  �          ����   $ %          � A � C       #  8'  �9   	   D       ��       ���� � �����  �  �          ����   ' (          � E � G       4  
(  P@      D       ��       ���� � �����  �  �          ����   ) *          � I � K       D  �(  �F      D       ��       ���� � �����  �  �          ����   + ,          � M � O       U  �)  pM      D       ��       ���� � �����  �  �          ����   - .          � Q � S       f  �*   T      D	       ��       ���� � �����  �  �          ����              � = � ?         �-  �      E        ��        ���� � �����  �  �          ����     !          � A � C       4  �.  x�      E       ��        ���� � �����  �  �          ����   " #          � E � G       J  �/  �      E       ��        ���� � �����  �  �          ����   $ %          � I � K       _  �0  X�   	   E       ��       ���� � �����  �  �          ����   & '          � M � O       u  �1  Ƚ      E       ��       ���� � �����  �  �          ����   ( )          � Q � S       �  x2  8�      E       ��       ���� � �����  �  �          ����   + ,          � U � W       �  h3  ��      E       ��       ���� � �����  �  �          ����   - .           Y  [       �  X4  �      E       ��       ���� � �����  �  �          ����   / 0          ] _       �  H5  ��      E       ��       ���� � �����  �  �          ����   1 2          a c       �  86  ��      E	       ��       ���� � -  �  �  �          ����   " #          � L � N       �  �9  �C      F      	  ��        ����	 � �����  �  �          ����   $ %          � P � R       �  ;  <N   
   F     	  ��        ����	 � �����  �  �          ����   & '          T V         <  �X      F     	  ��        ����	 � �����  �  �          ����   ( )          X Z         "=  Tc      F     	  ��       ����	 � �����  �  �          ����   * +          \ ^       8  0>  �m      F     	  ��       ����	 � �����  �  �          ����   , -          ` b       S  >?  lx      F     	  ��       ����	 � �����  �  �          ����   / 0          d f       n  L@  ��      F     	  ��       ����	 � �����  �  �          ����   1 2           h  j       �  ZA  ��      F     	  ��       ����	 � �����  �  �          ����   3 4          &l &n       �  hB  �       F     	  ��       ����	 � �����  �  �          ����   5 6          ,p ,r       �  vC  ��   ��  F	     	  ��       ����	 � 7  �  �  �           ����             � T - !       �   h  pb       �        ��        ���� � �������������          ����             � X 0 $         �  �e       �       ��        ���� � �������������          ����             � \ 3 '         �  xi       �       ��        ���� � �������������          ����             � ` 6 *         *  �l       �       ��       ���� � �������������          ����    !          � d 9 -          �  �p       �       ��       ���� � �������������          ����  " #          � h < 0       )  V  t       �       ��       ���� � �������������          ����  $ %          � l ? 3       2  �  �w       �       ��       ���� � �������������          ����  & '          � p B 6       ;  �  {       �       ��       ���� � �������������          ����  ) *          � t E 9       D    �~    
   �       ��       ���� � �������������          ����  + ,          � x H <       M  �  �    	   �	       ��       ���� � �������������           ����             � c 4 (       �    *�       �        ��        ���� � �������������          ����             � h 7 +       �  �  �       �       ��        ���� � �������������          ����    !          � m : .       �  n  �       �       ��        ���� � �������������          ����  # $          � r = 1       �  "  �       �       ��       ���� � �������������          ����  % &          � w @ 4       �  �  ڻ       �       ��       ���� � �������������          ����  ' (          � | C 7       �  �  ��       �       ��       ���� � �������������          ����  ) *          � � F :       �  >  ��       �       ��       ���� � �������������          ����  + ,          � � I =         �  ��    	   �       ��       ���� � �������������          ����  . /          � � L @         �  ��       �       ��       ���� � �������������          ����  0 1          � � O C         Z  v�       �	       ��       ���� � �������������          ����  ! "          � { : .       �  *!  P	      �        ��        ���� � �����  �  �          ����  # $          � � > 2       �  �!  �      �       ��        ���� � �����  �  �          ����  % &          � � B 6       �  �"  p      �       ��        ���� � �����  �  �          ����  ( )          � � F :       �  �#         �       ��       ���� � �����  �  �          ����  * +          � � J >       �  r$  �#      �       ��       ���� � �����  �  �          ����  , -          � � N B       �  D%   *   	   �       ��       ���� � �����  �  �          ����  . /          � � R F         &  �0      �       ��       ���� � �����  �  �          ����  0 1          � � V J         �&  @7      �       ��       ���� � �����  �  �          ����  3 4          � Z N       -  �'  �=      �       ��       ���� � �����  �  �          ����  5 6          
� ^ R       >  �(  `D      �	       ��       ���� � �����  �  �          ����  & '          � � J >       �  �+  t�      �        ��        ���� � �����  �  �          ����  ( )          � � N B         �,  �      �       ��        ���� � �����  �  �          ����  * +          � R F         �-  T�      �       ��        ���� � �����  �  �          ����  - .          	� V J       2  �.  ģ   	   �       ��       ���� � �����  �  �          ����  / 0          � Z N       H  �/  4�      �       ��       ���� � �����  �  �          ����  1 2          � ^ R       ]  �0  ��      �       ��       ���� � �����  �  �          ����  3 4          � b V       s  t1  �      �       ��       ���� � �����  �  �          ����  5 6          %� f Z       �  d2  ��      �       ��       ���� � �����  �  �          ����  8 9          ,� j ^       �  T3  ��      �       ��       ���� � �����  �  �          ����  : ;          3� n b       �  D4  d�      �	       ��       ���� � -  �  �  �          ����  + ,          � Y M       �  8  (0      �      	  ��        ����	 � �����  �  �          ����  - .          $� ] Q       �  9  �:   
   �     	  ��        ����	 � �����  �  �          ����  / 0          +� a U       �   :  @E      �     	  ��        ����	 � �����  �  �          ����  2 3          2� e Y       �  .;  �O      �     	  ��       ����	 � �����  �  �          ����  4 5          9� i ]         <<  XZ      �     	  ��       ����	 � �����  �  �          ����  6 7          @� m a       !  J=  �d      �     	  ��       ����	 � �����  �  �          ����  8 9          G� q e       <  X>  po      �     	  ��       ����	 � �����  �  �          ����  : ;          N� u i       W  f?  �y      �     	  ��       ����	 � �����  �  �          ����  = >          U� y m       r  t@  ��       �     	  ��       ����	 � �����  �  �          ����  ? @          \� } q       �  �A  �   ��  �	     	  ��       ����	 � 7  �  �  �           ����             , I � '       �   h  pb       �        ��        ���� � �������������          ����             / M � *         �  �e       �       ��        ���� � �������������          ����             2 Q � -         �  xi       �       ��        ���� � �������������          ����             5 U � 0         *  �l       �       ��       ���� � �������������          ����             8 Y � 3          �  �p       �       ��       ���� � �������������          ����             ; ] � 6       )  V  t       �       ��       ���� � �������������          ����              > a � 9       2  �  �w       �       ��       ���� � �������������          ����  ! "          A e � <       ;  �  {       �       ��       ���� � �������������          ����  # $          D i � ?       D    �~    
   �       ��       ���� � �������������          ����  % &          G m � B       M  �  �    	   �	       ��       ���� � �������������           ����             3 X � .       �    *�       �        ��        ���� � �������������          ����             7 \ � 1       �  �  �       �       ��        ���� � �������������          ����             ; ` � 4       �  n  �       �       ��        ���� � �������������          ����             ? d � 7       �  "  �       �       ��       ���� � �������������          ����             C h � :       �  �  ڻ       �       ��       ���� � �������������          ����  ! "          G l � =       �  �  ��       �       ��       ���� � �������������          ����  # $          K p � @       �  >  ��       �       ��       ���� � �������������          ����  % &          O t � C         �  ��    	   �       ��       ���� � �������������          ����  ' (          S x � F         �  ��       �       ��       ���� � �������������          ����  ) *          W | � I         Z  v�       �	       ��       ���� � �������������          ����             C g � 4       �  *!  P	      �        ��        ���� � �����  �  �          ����             G l � 8       �  �!  �      �       ��        ���� � �����  �  �          ����             K q � <       �  �"  p      �       ��        ���� � �����  �  �          ����    !          O v � @       �  �#         �       ��       ���� � �����  �  �          ����  " #          S { � D       �  r$  �#      �       ��       ���� � �����  �  �          ����  $ %          W � � H       �  D%   *   	   �       ��       ���� � �����  �  �          ����  ' (          [ � � L         &  �0      �       ��       ���� � �����  �  �          ����  ) *          _ � � P         �&  @7      �       ��       ���� � �����  �  �          ����  + ,          c � � T       -  �'  �=      �       ��       ���� � �����  �  �          ����  - .          g � X       >  �(  `D      �	       ��       ���� � �����  �  �          ����             S  � D       �  �+  t�      �        ��         ���� � �����  �  �          ����    !          W � � H         �,  �      �       ��         ���� � �����  �  �          ����  " #          [ � � L         �-  T�      �       ��         ���� � �����  �  �          ����  $ %          _ � P       2  �.  ģ   	   �       ��        ���� � �����  �  �          ����  & '          c � 	T       H  �/  4�      �       ��        ���� � �����  �  �          ����  ( )          g � X       ]  �0  ��      �       ��        ���� � �����  �  �          ����  + ,          k � \       s  t1  �      �       ��        ���� � �����  �  �          ����  - .          o � `       �  d2  ��      �       ��        ���� � �����  �  �          ����  / 0          s � %d       �  T3  ��      �       ��        ���� � �����  �  �          ����  1 2          w � ,h       �  D4  d�      �	       ��        ���� � -  �  �  �          ����  " #          b � S       �  8  (0      �      	  ��!        ����	 � �����  �  �          ����  $ %          f � W       �  9  �:   
   �     	  ��!        ����	 � �����  �  �          ����  & '          j � $[       �   :  @E      �     	  ��!        ����	 � �����  �  �          ����  ( )          n � +_       �  .;  �O      �     	  ��!       ����	 � �����  �  �          ����  * +          r � 2c         <<  XZ      �     	  ��!       ����	 � �����  �  �          ����  , -          v � 9g       !  J=  �d      �     	  ��!       ����	 � �����  �  �          ����  / 0          z � @k       <  X>  po      �     	  ��!       ����	 � �����  �  �          ����  1 2          ~ � Go       W  f?  �y      �     	  ��!       ����	 � �����  �  �          ����  3 4          � � Ns       r  t@  ��       �     	  ��!       ����	 � �����  �  �          ����  5 6          � � Uw       �  �A  �   ��  �	     	  ��!       ����	 � 7  �  �  �           ����                            ,  h       �        ��"        ���� � �������������           ����                            J  �       �       ��"        ���� � �������������           ����             !   !            h  �       �       ��"        ���� � �������������           ����             %   %            �         �       ��"       ���� � �������������           ����  	 
          )   )            �  H       �       ��"       ���� � �������������           ����             -   -         	   �  �       �       ��"       ���� � �������������           ����             1   1         	   �  �       �       ��"       ���� � �������������           ����             5   5         
   �  �       �       ��"       ���� � �������������           ����             9   9         
     8       �       ��"       ���� � �������������           ����             =   =            :  t       �	       ��"       ���� � �������������           ����             +  +            �         �        ��#        ���� � �������������           ����             /  /            �  �       �       ��#        ���� � �������������           ����  	 
          3  3            *  ~	       �       ��#        ���� � �������������           ����             7  7            f  2
       �       ��#       ���� � �������������           ����             ;  ;            �  �
       �       ��#       ���� � �������������           ����             ?  ?            �  �       �       ��#       ���� � �������������           ����             C  C              N       �       ��#       ���� � �������������           ����             G ! G         !   V         �       ��#       ���� � �������������           ����             K # K         #   �  �       �       ��#       ���� � �������������           ����             O % O         $   �  j       �	       ��#       ���� � �������������           ����  	 
          <  <        :   �  �       �        ��$        ���� � �������������          ����             A  A        >     `       �       ��$        ���� � �������������          ����             F  F        B   r  �       �       ��$        ���� � �������������          ����             K  K        E   �  0       �       ��$       ���� � �������������          ����             P  P        I   &  �       �       ��$       ���� � �������������          ����             U   U "       L   �          �       ��$       ���� � �������������          ����             Z # Z %       P   �  h       �       ��$       ���� � �������������          ����             _ & _ (       T   4  �        �       ��$       ���� � �������������          ����             d ) d +       W   �  8"       �       ��$       ���� � �������������          ����             i , i .       [   �  �#       �	       ��$       ���� � �������������           ����             V  V        �   P
  �3       �        ��%        ���� � �������������          ����             [  [        �   �
  �5       �       ��%        ���� � �������������          ����             `  ` !       �   @  @8       �       ��%        ���� � �������������          ����             e " e $       �   �  �:       �       ��%       ���� � �������������          ����             j % j '       �   0  �<       �       ��%       ���� � �������������          ����             o ( o *       �   �  H?       �       ��%       ���� � �������������          ����             t + t -       �      �A       �       ��%       ���� � �������������          ����             y . y 0       �   �  �C       �       ��%       ���� � �������������          ����             ~ 1 ~ 3       �     PF       �       ��%       ���� � �������������          ����    !          � 4 � 6       �   �  �H       �	       ��%       ���� � �������������           ����             o   o "       �   h  pb       �        ��&        ���� � �������������          ����             t # t %         �  �e       �       ��&        ���� � �������������          ����             y & y (         �  xi       �       ��&        ���� � �������������          ����             ~ ) ~ +         *  �l       �       ��&       ���� � �������������          ����             � , � .          �  �p       �       ��&       ���� � �������������          ����             � / � 1       )  V  t       �       ��&       ���� � �������������          ����             � 2 � 4       2  �  �w       �       ��&       ���� � �������������          ����    !          � 5 � 7       ;  �  {       �       ��&       ���� � �������������          ����  " #          � 8 � :       D    �~    
   �       ��&       ���� � �������������          ����  $ %          � ; � =       M  �  �    	   �	       ��&       ���� � �������������           ����             � ' � )       �    *�       �        ��'        ���� � �������������          ����             � * � ,       �  �  �       �       ��'        ���� � �������������          ����             � - � /       �  n  �       �       ��'        ���� � �������������          ����             � 0 � 2       �  "  �       �       ��'       ���� � �������������          ����             � 3 � 5       �  �  ڻ       �       ��'       ���� � �������������          ����    !          � 6 � 8       �  �  ��       �       ��'       ���� � �������������          ����  " #          � 9 � ;       �  >  ��       �       ��'       ���� � �������������          ����  $ %          � < � >         �  ��    	   �       ��'       ���� � �������������          ����  & '          � ? � A         �  ��       �       ��'       ���� � �������������          ����  ( )          � B � D         Z  v�       �	       ��'       ���� � �������������          ����             � - � /       �  *!  P	      �        ��(        ���� � �����  �  �          ����             � 1 � 3       �  �!  �      �       ��(        ���� � �����  �  �          ����             � 5 � 7       �  �"  p      �       ��(        ���� � �����  �  �          ����              � 9 � ;       �  �#         �       ��(       ���� � �����  �  �          ����  ! "          � = � ?       �  r$  �#      �       ��(       ���� � �����  �  �          ����  $ %          � A � C       �  D%   *   	   �       ��(       ���� � �����  �  �          ����  & '          � E � G         &  �0      �       ��(       ���� � �����  �  �          ����  ( )          � I � K         �&  @7      �       ��(       ���� � �����  �  �          ����  * +          � M � O       -  �'  �=      �       ��(       ���� � �����  �  �          ����  , -          � Q � S       >  �(  `D      �	       ��(       ���� � �����  �  �          ����             � = � ?       �  �+  t�      �        ��)        ���� � �����  �  �          ����              � A � C         �,  �      �       ��)        ���� � �����  �  �          ����  ! "          � E � G         �-  T�      �       ��)        ���� � �����  �  �          ����  # $          � I � K       2  �.  ģ   	   �       ��)       ���� � �����  �  �          ����  % &          � M � O       H  �/  4�      �       ��)       ���� � �����  �  �          ����  ' (          � Q � S       ]  �0  ��      �       ��)       ���� � �����  �  �          ����  * +          � U � W       s  t1  �      �       ��)       ���� � �����  �  �          ����  , -          � Y � [       �  d2  ��      �       ��)       ���� � �����  �  �          ����  . /          � ] � _       �  T3  ��      �       ��)       ���� � �����  �  �          ����  0 1          � a � c       �  D4  d�      �	       ��)       ���� � -  �  �  �          ����  ! "          � L � N       �  8  (0      �      	  ��*        ����	 � �����  �  �          ����  # $          � P � R       �  9  �:   
   �     	  ��*        ����	 � �����  �  �          ����  % &          � T � V       �   :  @E      �     	  ��*        ����	 � �����  �  �          ����  ' (          � X � Z       �  .;  �O      �     	  ��*       ����	 � �����  �  �          ����  ) *          � \ � ^         <<  XZ      �     	  ��*       ����	 � �����  �  �          ����  + ,          � ` � b       !  J=  �d      �     	  ��*       ����	 � �����  �  �          ����  . /          d f       <  X>  po      �     	  ��*       ����	 � �����  �  �          ����  0 1          h j       W  f?  �y      �     	  ��*       ����	 � �����  �  �          ����  2 3          l n       r  t@  ��       �     	  ��*       ����	 � �����  �  �          ����  4 5          p r       �  �A  �   ��  �	     	  ��*       ����	 � 7  �  �  �          
 ��              � T - ! F     ����,  �        �       �    +        ���� � �������������          
 ��              � X 0 $ F     �����  ��        �      �    +        ���� � �������������          
 ��              � \ 3 ' F     ����X  �        �      �    +        ���� � �������������           ��  ! "           � ` 6 * F     �����  ��        �      �    +        ���� � �������������           ��  # $           � d 9 - F     �����  �        �      �    +        ���� � �������������           ��  % &           � h < 0 F     ����  ��        �      �    +        ���� � �������������           ��  ' (           � l ? 3 F     �����   �        �      �    +        ���� � �������������           ��  ) *           � p B 6 F     ����F  ��        �      �    +        ���� � �������������           ��  , -           � t E 9 F     �����  (�        �      �    +        ���� � �������������           ��  . /           � x H < F     ����r  ��        � 	     �    +        ���� � �������������           ��               � c 4 ( P     �����!  ��        �       �    ,        ���� � �������������           ��  ! "           � h 7 + P     ����~"  r�        �      �    ,        ���� � �������������           ��  # $           � m : . P     ����2#  ^�        �      �    ,        ���� � �������������           ��  & '           � r = 1 P     �����#  J�        �      �    ,        ���� � �������������           ��  ( )           � w @ 4 P     �����$  6        �      �    ,        ���� � �������������           ��  * +           � | C 7 P     ����N%  "       �      �    ,        ���� � �������������           ��  , -           � � F : P     ����&  
       �      �    ,        ���� � �������������           ��  . /           � I = P     �����&  �       �      �    ,        ���� � �������������           ��  1 2           
� L @ P     ����j'  �       �      �    ,        ���� � �������������           ��  3 4           � O C P     ����(  �       � 	     �    ,        ���� � �������������           ��  $ %           � { : . Z     �����*  pW       �       �    -        ���� � �����  �  �           ��  & '           � > 2 Z     �����+   ^       �      �    -        ���� � �����  �  �           ��  ( )           � B 6 Z     �����,  �d       �      �    -        ���� � �����  �  �           ��  + ,           � F : Z     ����d-   k       �      �    -        ���� � �����  �  �           ��  - .           � J > Z     ����6.  �q       �      �    -        ���� � �����  �  �           ��  / 0           � N B Z     ����/  @x       �      �    -        ���� � �����  �  �           ��  1 2           � R F Z     �����/  �~       �      �    -        ���� � �����  �  �           ��  3 4           %� V J Z     �����0  `�       �      �    -        ���� � �����  �  �           ��  6 7           +� Z N Z     ����~1  ��       �      �    -        ���� � �����  �  �           ��  8 9           1� ^ R Z     ����P2  ��       � 	     �    -        ���� � �����  �  �           ��  ) *           � J > d     �����5  X�       �       �    .        ���� � �����  �  �           ��  + ,           "� N B d     �����6  ��       �      �    .        ���� � �����  �  �           ��  - .           )� R F d     ����x7  8�       �      �    .        ���� � �����  �  �           ��  0 1           0� V J d     ����h8  ��       �      �    .        ���� � �����  �  �           ��  2 3           7� Z N d     ����X9         �      �    .        ���� � �����  �  �           ��  4 5           >� ^ R d     ����H:  �       �      �    .        ���� � �����  �  �           ��  6 7           E� b V d     ����8;  �       �      �    .        ���� � �����  �  �           ��  8 9           L� f Z d     ����(<  h       �      �    .        ���� � �����  �  �           ��  ; <           S� j ^ d     ����=  �%       �      �    .        ���� � �����  �  �           ��  = >           Z� n b d     ����>  H.       � 	     �    .        ���� � �����  �  �           ��  . /           D� Y M n     �����A  Б       �       �    /        ����	 � �����  �  �           ��  0 1           K� ] Q n     �����B  \�       �      �    /        ����	 � �����  �  �           ��  2 3           R� a U n     �����C  �       �      �    /        ����	 � �����  �  �           ��  5 6           Y� e Y n     �����D  t�       �      �    /        ����	 � �����  �  �           ��  7 8           `� i ] n     ���� F   �       �      �    /        ����	 � �����  �  �           ��  9 :           g� m a n     ����G  ��       �      �    /        ����	 � �����  �  �           ��  ; <           n� q e n     ����H  �       �      �    /        ����	 � �����  �  �           ��  = >           u� u i n     ����*I  ��       �      �    /        ����	 � �����  �  �           ��  @ A           |� y m n     ����8J  0�       �      �    /        ����	 � �����  �  �           ��  B C           �� } q n     ����FK  ��       � 	     �    /        ����	 � �����  �  �          
 ��              R p � ' F     ����,  �        �       �    0        ���� � �������������          
 ��              U t � * F     �����  ��        �      �    0        ���� � �������������          
 ��              X x � - F     ����X  �        �      �    0        ���� � �������������           ��              [ | � 0 F     �����  ��        �      �    0        ���� � �������������           ��              ^ � � 3 F     �����  �        �      �    0        ���� � �������������           ��              a � � 6 F     ����  ��        �      �    0        ���� � �������������           ��    !           d � � 9 F     �����   �        �      �    0        ���� � �������������           ��  " #           g � � < F     ����F  ��        �      �    0        ���� � �������������           ��  $ %           j � � ? F     �����  (�        �      �    0        ���� � �������������           ��  & '           m � � B F     ����r  ��        � 	     �    0        ���� � �������������           ��              Y  � . P     �����!  ��        �       �    1        ���� � �������������           ��              ] � � 1 P     ����~"  r�        �      �    1        ���� � �������������           ��              a � � 4 P     ����2#  ^�        �      �    1        ���� � �������������           ��              e � � 7 P     �����#  J�        �      �    1        ���� � �������������           ��               i � � : P     �����$  6        �      �    1        ���� � �������������           ��  " #           m � � = P     ����N%  "       �      �    1        ���� � �������������           ��  $ %           q � � @ P     ����&  
       �      �    1        ���� � �������������           ��  & '           u � � C P     �����&  �       �      �    1        ���� � �������������           ��  ( )           y � F P     ����j'  �       �      �    1        ���� � �������������           ��  * +           } � 	I P     ����(  �       � 	     �    1        ���� � �������������           ��              i � � 4 Z     �����*  pW       �       �    2        ���� � �����  �  �           ��              m � � 8 Z     �����+   ^       �      �    2        ���� � �����  �  �           ��               q �  < Z     �����,  �d       �      �    2        ���� � �����  �  �           ��  ! "           u � @ Z     ����d-   k       �      �    2        ���� � �����  �  �           ��  # $           y � D Z     ����6.  �q       �      �    2        ���� � �����  �  �           ��  % &           } � H Z     ����/  @x       �      �    2        ���� � �����  �  �           ��  ( )           � � L Z     �����/  �~       �      �    2        ���� � �����  �  �           ��  * +           � � P Z     �����0  `�       �      �    2        ���� � �����  �  �           ��  , -           � � $T Z     ����~1  ��       �      �    2        ���� � �����  �  �           ��  . /           � � *X Z     ����P2  ��       � 	     �    2        ���� � �����  �  �           ��               y � D d     �����5  X�       �       �    3        ���� � �����  �  �           ��  ! "           } � H d     �����6  ��       �      �    3        ���� � �����  �  �           ��  # $           � � "L d     ����x7  8�       �      �    3        ���� � �����  �  �           ��  % &           � � )P d     ����h8  ��       �      �    3        ���� � �����  �  �           ��  ' (           � � 0T d     ����X9         �      �    3        ���� � �����  �  �           ��  ) *           � � 7X d     ����H:  �       �      �    3        ���� � �����  �  �           ��  , -           � � >\ d     ����8;  �       �      �    3        ���� � �����  �  �           ��  . /           � � E` d     ����(<  h       �      �    3        ���� � �����  �  �           ��  0 1           � � Ld d     ����=  �%       �      �    3        ���� � �����  �  �           ��  2 3           � � Sh d     ����>  H.       � 	     �    3        ���� � �����  �  �           ��  # $           � � =S n     �����A  Б       �       �    4        ����	 � �����  �             ��  % &           � � DW n     �����B  \�       �      �    4        ����	 � �����  �             ��  ' (           � � K[ n     �����C  �       �      �    4        ����	 � �����  �             ��  ) *           � � R_ n     �����D  t�       �      �    4        ����	 � �����  �             ��  + ,           � � Yc n     ���� F   �       �      �    4        ����	 � �����  �             ��  - .           � � `g n     ����G  ��       �      �    4        ����	 � �����  �             ��  0 1           � � gk n     ����H  �       �      �    4        ����	 � �����  �             ��  2 3           � � no n     ����*I  ��       �      �    4        ����	 � �����  �             ��  4 5           � � us n     ����8J  0�       �      �    4        ����	 � �����  �             ��  6 7           � � |w n     ����FK  ��       � 	     �    4        ����	 � �����  �               ��              @   @        �����
  �         �       �    5        ���� � ������������            ��              D   D        ����          �      �    5        ���� � ������������            ��              H   H        ����,  X        �      �    5        ���� � ������������            ��   	           L   L        ����J  �        �      �    5        ���� � ������������            ��  
            P   P        ����h  �        �      �    5        ���� � ������������            ��              T   T        �����          �      �    5        ���� � ������������            ��              X   X        �����  H        �      �    5        ���� � ������������            ��              \   \        �����  �        �      �    5        ���� � ������������            ��              `   `        �����  �        �      �    5        ���� � ������������            ��              d   d        �����  �        � 	     �    5        ���� � ������������           ��              R  R   (     ����v  b%        �       �    6        ���� � ������������           ��   	           V  V   (     �����  &        �      �    6        ���� � ������������           ��  
            Z  Z   (     �����  �&        �      �    6        ���� � ������������           ��              ^  ^   (     ����*  ~'        �      �    6        ���� � ������������           ��              b  b   (     ����f  2(        �      �    6        ���� � ������������           ��              f  f   (     �����  �(        �      �    6        ���� � ������������           ��              j  j   (     �����  �)        �      �    6        ���� � ������������           ��              n ! n   (     ����  N*        �      �    6        ���� � ������������           ��              r # r   (     ����V  +        �      �    6        ���� � ������������           ��              v % v   (     �����  �+        � 	     �    6        ���� � ������������          ��  
            c  c  2     �����  >        �       �    7        ���� � ������������          ��              h  h  2     �����  p?        �      �    7        ���� � ������������          ��              m  m  2     ����6  �@        �      �    7        ���� � ������������          ��              r  r  2     �����  @B        �      �    7        ���� � ������������          ��              w  w  2     �����  �C        �      �    7        ���� � ������������          ��              |   | " 2     ����D  E        �      �    7        ���� � ������������          ��              � # � % 2     �����  xF        �      �    7        ���� � ������������          ��              � & � ( 2     �����  �G        �      �    7        ���� � ������������          ��              � ) � + 2     ����R  HI        �      �    7        ���� � ������������          ��              � , � . 2     �����  �J        � 	     �    7        ���� � ������������         	 ��              }  }  <     ����  dd        �       �    8        ���� � ������������         	 ��              �  �  <     �����  �f        �      �    8        ���� � ������������         	 ��              �  � ! <     ����  i        �      �    8        ���� � ������������         	 ��              � " � $ <     ����|  lk        �      �    8        ���� � ������������         	 ��              � % � ' <     �����  �m        �      �    8        ���� � ������������         	 ��              � ( � * <     ����l  p        �      �    8        ���� � ������������         	 ��              � + � - <     �����  tr        �      �    8        ���� � ������������         	 ��              � . � 0 <     ����\  �t        �      �    8        ���� � ������������         	 ��               � 1 � 3 <     �����  $w        �      �    8        ���� � ������������         	 ��  ! "           � 4 � 6 <     ����L  |y        � 	     �    8        ���� � ������������         
 ��              �   � " F     ����,  �        �       �    9        ���� � ������������         
 ��              � # � % F     �����  ��        �      �    9        ���� � ������������         
 ��              � & � ( F     ����X  �        �      �    9        ���� � ������������          ��              � ) � + F     �����  ��        �      �    9        ���� � ������������          ��              � , � . F     �����  �        �      �    9        ���� � ������������          ��              � / � 1 F     ����  ��        �      �    9        ���� � ������������          ��               � 2 � 4 F     �����   �        �      �    9        ���� � ������������          ��  ! "           � 5 � 7 F     ����F  ��        �      �    9        ���� � ������������          ��  # $           � 8 � : F     �����  (�        �      �    9        ���� � ������������          ��  % &           � ; � = F     ����r  ��        � 	     �    9        ���� � ������������          ��              � ' � ) P     �����!  ��        �       �    :        ���� � ������������          ��              � * � , P     ����~"  r�        �      �    :        ���� � ������������          ��              � - � / P     ����2#  ^�        �      �    :        ���� � ������������          ��              � 0 � 2 P     �����#  J�        �      �    :        ���� � ������������          ��              � 3 � 5 P     �����$  6        �      �    :        ���� � ������������          ��  ! "           � 6 � 8 P     ����N%  "       �      �    :        ���� � ������������          ��  # $           � 9 � ; P     ����&  
       �      �    :        ���� � ������������          ��  % &           � < � > P     �����&  �       �      �    :        ���� � ������������          ��  ' (           � ? � A P     ����j'  �       �      �    :        ���� � ������������          ��  ) *           � B � D P     ����(  �       � 	     �    :        ���� � ������������          ��              � - � / Z     �����*  pW       �       �    ;        ���� � �����  �            ��              � 1 � 3 Z     �����+   ^       �      �    ;        ���� � �����  �            ��              � 5 � 7 Z     �����,  �d       �      �    ;        ���� � �����  �            ��    !           � 9 � ; Z     ����d-   k       �      �    ;        ���� � �����  �            ��  " #           � = � ? Z     ����6.  �q       �      �    ;        ���� � �����  �            ��  $ %           � A � C Z     ����/  @x       �      �    ;        ���� � �����  �            ��  ' (           � E � G Z     �����/  �~       �      �    ;        ���� � �����  �            ��  ) *           � I � K Z     �����0  `�       �      �    ;        ���� � �����  �            ��  + ,           � M � O Z     ����~1  ��       �      �    ;        ���� � �����  �            ��  - .           � Q � S Z     ����P2  ��       � 	     �    ;        ���� � �����  �            ��              � = � ? d     �����5  X�       �       �    <        ���� � �����  �            ��    !           � A � C d     �����6  ��       �      �    <        ���� � �����  �            ��  " #           � E � G d     ����x7  8�       �      �    <        ���� � �����  �            ��  $ %           � I � K d     ����h8  ��       �      �    <        ���� � �����  �            ��  & '            M  O d     ����X9         �      �    <        ���� � �����  �            ��  ( )           Q S d     ����H:  �       �      �    <        ���� � �����  �            ��  + ,           U W d     ����8;  �       �      �    <        ���� � �����  �            ��  - .           Y [ d     ����(<  h       �      �    <        ���� � �����  �            ��  / 0           ] _ d     ����=  �%       �      �    <        ���� � �����  �            ��  1 2           a c d     ����>  H.       � 	     �    <        ���� � �����  �            ��  " #           L N n     �����A  Б       �       �    =        ����	 � �����  �  	          ��  $ %           P R n     �����B  \�       �      �    =        ����	 � �����  �  	          ��  & '           T V n     �����C  �       �      �    =        ����	 � �����  �  	          ��  ( )           X Z n     �����D  t�       �      �    =        ����	 � �����  �  	          ��  * +            \  ^ n     ���� F   �       �      �    =        ����	 � �����  �  	          ��  , -           &` &b n     ����G  ��       �      �    =        ����	 � �����  �  	          ��  / 0           ,d ,f n     ����H  �       �      �    =        ����	 � �����  �  	          ��  1 2           2h 2j n     ����*I  ��       �      �    =        ����	 � �����  �  	          ��  3 4           8l 8n n     ����8J  0�       �      �    =        ����	 � �����  �  	          ��  5 6           >p >r n     ����FK  ��       � 	     �    =        ����	 � �����  �  	         ����             � T - !       �     `       �        ��>        ���� � ������������
         ����             � X 0 $       �   �  �c       �       ��>        ���� � ������������
         ����             � \ 3 '         0   g       �       ��>        ���� � ������������
         ����              � ` 6 *         �  �j       �       ��>       ���� � ������������
         ����  ! "          � d 9 -         \  (n       �       ��>       ���� � ������������
         ����  # $          � h < 0       #  �  �q       �       ��>       ���� � ������������
         ����  % &          � l ? 3       ,  �  0u       �       ��>       ���� � ������������
         ����  ' (          � p B 6       5    �x       �       ��>       ���� � ������������
         ����  * +          � t E 9       >  �  8|    
   �       ��>       ���� � ������������
         ����  , -          � x H <       G  J  �    	   �	       ��>       ���� � ������������
         ����             � c 4 (       �  �  n�       �        ��?        ���� � ������������         ����              � h 7 +       �  V  Z�       �       ��?        ���� � ������������         ����  ! "          � m : .       �  
  F�       �       ��?        ���� � ������������         ����  $ %          � r = 1       �  �  2�       �       ��?       ���� � ������������         ����  & '          � w @ 4       �  r  �       �       ��?       ���� � ������������         ����  ( )          � | C 7       �  &  
�       �       ��?       ���� � ������������         ����  * +          � � F :       �  �  ��       �       ��?       ���� � ������������         ����  , -          � � I =       �  �  ��    	   �       ��?       ���� � ������������         ����  / 0          � � L @         B  ��       �       ��?       ���� � ������������         ����  1 2          � � O C         �  ��       �	       ��?       ���� � ������������         ����  " #          � { : .       �  �   0      �        ��@        ���� � �����  �           ����  $ %          � � > 2       �  �!  �      �       ��@        ���� � �����  �           ����  & '          � � B 6       �  j"  P      �       ��@        ���� � �����  �           ����  ) *          � � F :       �  <#  �      �       ��@       ���� � �����  �           ����  + ,          � � J >       �  $  p       �       ��@       ���� � �����  �           ����  - .          � � N B       �  �$   '   	   �       ��@       ���� � �����  �           ����  / 0          � R F         �%  �-      �       ��@       ���� � �����  �           ����  1 2          � V J         �&   4      �       ��@       ���� � �����  �           ����  4 5          � Z N       %  V'  �:      �       ��@       ���� � �����  �           ����  6 7          � ^ R       6  ((  @A      �	       ��@       ���� � �����  �           ����  ' (          � J >       �  p+  ��      �        ��A        ���� � �����  �           ����  ) *          � N B       �  `,  `�      �       ��A        ���� � �����  �           ����  + ,          � R F         P-  З      �       ��A        ���� � �����  �           ����  . /          � V J       )  @.  @�   	   �       ��A       ���� � �����  �           ����  0 1          � Z N       ?  0/  ��      �       ��A       ���� � �����  �           ����  2 3          $� ^ R       T   0   �      �       ��A       ���� � �����  �           ����  4 5          +� b V       j  1  ��      �       ��A       ���� � �����  �           ����  6 7          2� f Z       �   2   �      �       ��A       ���� � �����  �           ����  9 :          9� j ^       �  �2  p�      �       ��A       ���� � �����  �           ����  ; <          @� n b       �  �3  ��      �	       ��A       ���� � -  �  �           ����  , -          *� Y M       �  �7  @,      �      	  ��B        ����	 � �����  �           ����  . /          1� ] Q       �  �8  �6   
   �     	  ��B        ����	 � �����  �           ����  0 1          8� a U       �  �9  XA      �     	  ��B        ����	 � �����  �           ����  3 4          ?� e Y       �  �:  �K      �     	  ��B       ����	 � �����  �           ����  5 6          F� i ]       �  �;  pV      �     	  ��B       ����	 � �����  �           ����  7 8          M� m a         �<  �`      �     	  ��B       ����	 � �����  �           ����  9 :          T� q e       2  �=  �k      �     	  ��B       ����	 � �����  �           ����  ; <          [� u i       M  ?  v      �     	  ��B       ����	 � �����  �           ����  > ?          b� y m       h  @  ��       �     	  ��B       ����	 � �����  �           ����  @ A          i� } q       �  A  ,�   ��  �	     	  ��B       ����	 � 7  �  �           ����             9 V � '       �     `               ��C        ���� � ������������         ����             < Z � *       �   �  �c              ��C        ���� � ������������         ����             ? ^ � -         0   g              ��C        ���� � ������������         ����             B b � 0         �  �j              ��C       ���� � ������������         ����             E f � 3         \  (n              ��C       ���� � ������������         ����             H j � 6       #  �  �q              ��C       ���� � ������������         ����              K n � 9       ,  �  0u              ��C       ���� � ������������         ����  ! "          N r � <       5    �x              ��C       ���� � ������������         ����  # $          Q v � ?       >  �  8|    
          ��C       ���� � ������������         ����  % &          T z � B       G  J  �    	   	       ��C       ���� � ������������         ����             @ e � .       �  �  n�               ��D        ���� � ������������         ����             D i � 1       �  V  Z�              ��D        ���� � ������������         ����             H m � 4       �  
  F�              ��D        ���� � ������������         ����             L q � 7       �  �  2�              ��D       ���� � ������������         ����             P u � :       �  r  �              ��D       ���� � ������������         ����  ! "          T y � =       �  &  
�              ��D       ���� � ������������         ����  # $          X } � @       �  �  ��              ��D       ���� � ������������         ����  % &          \ � � C       �  �  ��    	          ��D       ���� � ������������         ����  ' (          ` � � F         B  ��              ��D       ���� � ������������         ����  ) *          d � � I         �  ��       	       ��D       ���� � ������������         ����             P t � 4       �  �   0              ��E        ���� � �����  �           ����             T y � 8       �  �!  �             ��E        ���� � �����  �           ����             X ~ � <       �  j"  P             ��E        ���� � �����  �           ����    !          \ � � @       �  <#  �             ��E       ���� � �����  �           ����  " #          ` � � D       �  $  p              ��E       ���� � �����  �           ����  $ %          d � � H       �  �$   '   	          ��E       ���� � �����  �           ����  ' (          h � � L         �%  �-             ��E       ���� � �����  �           ����  ) *          l � P         �&   4             ��E       ���� � �����  �           ����  + ,          p � 
T       %  V'  �:             ��E       ���� � �����  �           ����  - .          t � X       6  ((  @A      	       ��E       ���� � �����  �           ����             ` � � D       �  p+  ��              ��F        ���� � �����  �           ����    !          d � H       �  `,  `�             ��F        ���� � �����  �           ����  " #          h � L         P-  З             ��F        ���� � �����  �           ����  $ %          l � P       )  @.  @�   	          ��F       ���� � �����  �           ����  & '          p � T       ?  0/  ��             ��F       ���� � �����  �           ����  ( )          t � X       T   0   �             ��F       ���� � �����  �           ����  + ,          x � $\       j  1  ��             ��F       ���� � �����  �           ����  - .          | � +`       �   2   �             ��F       ���� � �����  �           ����  / 0          � � 2d       �  �2  p�             ��F       ���� � �����  �           ����  1 2          � � 9h       �  �3  ��      	       ��F       ���� � -  �  �           ����  " #          o � #S       �  �7  @,      	      	  ��G        ����	 � �����  �           ����  $ %          s � *W       �  �8  �6   
   	     	  ��G        ����	 � �����  �           ����  & '          w � 1[       �  �9  XA      	     	  ��G        ����	 � �����  �           ����  ( )          { � 8_       �  �:  �K      	     	  ��G       ����	 � �����  �           ����  * +           � ?c       �  �;  pV      	     	  ��G       ����	 � �����  �           ����  , -          � � Fg         �<  �`      	     	  ��G       ����	 � �����  �           ����  / 0          � � Mk       2  �=  �k      	     	  ��G       ����	 � �����  �           ����  1 2          � � To       M  ?  v      	     	  ��G       ����	 � �����  �           ����  3 4          � � [s       h  @  ��       	     	  ��G       ����	 � �����  �           ����  5 6          � � bw       �  A  ,�   ��  		     	  ��G       ����	 � 7  �  �            ����             &   &            �   �                ��H        ���� � ������������          ����             *   *            �   �              ��H        ���� � ������������          ����             .   .                            ��H        ���� � ������������          ����             2   2            "  D              ��H       ���� � ������������          ����  	 
          6   6            @  �              ��H       ���� � ������������          ����             :   :            ^  �              ��H       ���� � ������������          ����             >   >            |  �              ��H       ���� � ������������          ����             B   B            �  4              ��H       ���� � ������������          ����             F   F            �  p              ��H       ���� � ������������          ����             J   J         	   �  �       	       ��H       ���� � ������������          ����             8  8            N  �               ��I        ���� � ������������          ����             <  <            �  �              ��I        ���� � ������������          ����  	 
          @  @            �  R              ��I        ���� � ������������          ����             D  D              	              ��I       ���� � ������������          ����             H  H            >  �	              ��I       ���� � ������������          ����             L  L            z  n
              ��I       ���� � ������������          ����             P  P            �  "              ��I       ���� � ������������          ����             T ! T            �  �              ��I       ���� � ������������          ����             X # X             .  �              ��I       ���� � ������������          ����             \ % \         !   j  >       	       ��I       ���� � ������������         ����  	 
          I  I        6   Z  h               ��J        ���� � ������������         ����             N  N        :   �  �              ��J        ���� � ������������         ����             S  S        >     8              ��J        ���� � ������������         ����             X  X        A   h  �              ��J       ���� � ������������         ����             ]  ]        E   �                ��J       ���� � ������������         ����             b   b "       H     p              ��J       ���� � ������������         ����             g # g %       L   v  �              ��J       ���� � ������������         ����             l & l (       P   �  @              ��J       ���� � ������������         ����             q ) q +       S   *  �               ��J       ���� � ������������         ����             v , v .       W   �  "       	       ��J       ���� � ������������         ����             c  c           �	  �1               ��K        ���� � ������������         ����             h  h        �   d
  �3              ��K        ���� � ������������         ����             m  m !       �   �
  L6              ��K        ���� � ������������         ����             r " r $       �   T  �8              ��K       ���� � ������������         ����             w % w '       �   �  �:              ��K       ���� � ������������         ����             | ( | *       �   D  T=              ��K       ���� � ������������         ����             � + � -       �   �  �?              ��K       ���� � ������������         ����             � . � 0       �   4  B              ��K       ���� � ������������         ����             � 1 � 3       �   �  \D              ��K       ���� � ������������         ����    !          � 4 � 6       �   $  �F       	       ��K       ���� � ������������         ����             |   | "       �     `               ��L        ���� � ������������         ����             � # � %       �   �  �c              ��L        ���� � ������������         ����             � & � (         0   g              ��L        ���� � ������������         ����             � ) � +         �  �j              ��L       ���� � ������������         ����             � , � .         \  (n              ��L       ���� � ������������         ����             � / � 1       #  �  �q              ��L       ���� � ������������         ����             � 2 � 4       ,  �  0u              ��L       ���� � ������������         ����    !          � 5 � 7       5    �x              ��L       ���� � ������������         ����  " #          � 8 � :       >  �  8|    
          ��L       ���� � ������������         ����  $ %          � ; � =       G  J  �    	   	       ��L       ���� � ������������         ����             � ' � )       �  �  n�               ��M        ���� � ������������         ����             � * � ,       �  V  Z�              ��M        ���� � ������������         ����             � - � /       �  
  F�              ��M        ���� � ������������         ����             � 0 � 2       �  �  2�              ��M       ���� � ������������         ����             � 3 � 5       �  r  �              ��M       ���� � ������������         ����    !          � 6 � 8       �  &  
�              ��M       ���� � ������������         ����  " #          � 9 � ;       �  �  ��              ��M       ���� � ������������         ����  $ %          � < � >       �  �  ��    	          ��M       ���� � ������������         ����  & '          � ? � A         B  ��              ��M       ���� � ������������         ����  ( )          � B � D         �  ��       	       ��M       ���� � ������������         ����             � - � /       �  �   0              ��N        ���� � �����  �           ����             � 1 � 3       �  �!  �             ��N        ���� � �����  �           ����             � 5 � 7       �  j"  P             ��N        ���� � �����  �           ����              � 9 � ;       �  <#  �             ��N       ���� � �����  �           ����  ! "          � = � ?       �  $  p              ��N       ���� � �����  �           ����  $ %          � A � C       �  �$   '   	          ��N       ���� � �����  �           ����  & '          � E � G         �%  �-             ��N       ���� � �����  �           ����  ( )          � I � K         �&   4             ��N       ���� � �����  �           ����  * +          � M � O       %  V'  �:             ��N       ���� � �����  �           ����  , -          � Q � S       6  ((  @A      	       ��N       ���� � �����  �           ����             � = � ?       �  p+  ��              ��O        ���� � �����  �           ����              � A � C       �  `,  `�             ��O        ���� � �����  �           ����  ! "          � E � G         P-  З             ��O        ���� � �����  �           ����  # $          � I � K       )  @.  @�   	          ��O       ���� � �����  �           ����  % &          � M � O       ?  0/  ��             ��O       ���� � �����  �           ����  ' (          � Q � S       T   0   �             ��O       ���� � �����  �           ����  * +          � U � W       j  1  ��             ��O       ���� � �����  �           ����  , -          � Y � [       �   2   �             ��O       ���� � �����  �           ����  . /          � ] � _       �  �2  p�             ��O       ���� � �����  �           ����  0 1          a c       �  �3  ��      	       ��O       ���� � -  �  �           ����  ! "          � L � N       �  �7  @,            	  ��P        ����	 � �����  �           ����  # $          � P � R       �  �8  �6   
        	  ��P        ����	 � �����  �           ����  % &          � T � V       �  �9  XA           	  ��P        ����	 � �����  �           ����  ' (           X  Z       �  �:  �K           	  ��P       ����	 � �����  �           ����  ) *          \ ^       �  �;  pV           	  ��P       ����	 � �����  �           ����  + ,          ` b         �<  �`           	  ��P       ����	 � �����  �           ����  . /          d f       2  �=  �k           	  ��P       ����	 � �����  �           ����  0 1          h j       M  ?  v           	  ��P       ����	 � �����  �           ����  2 3          l n       h  @  ��            	  ��P       ����	 � �����  �           ����  4 5          $p $r       �  A  ,�   ��  	     	  ��P       ����	 � 7  �  �            ����             � T - !       b    H�       Z        ��Q        ���� � ������������         ����             � X 0 $       k  �  ̍       Z       ��Q        ���� � ������������         ����             � \ 3 '       t  8  P�       Z       ��Q        ���� � ������������         ����             � ` 6 *       }  �  Ԕ       Z       ��Q       ���� � ������������         ����    !          � d 9 -       �  d  X�       Z       ��Q       ���� � ������������         ����  " #          � h < 0       �  �  ܛ       Z       ��Q       ���� � ������������         ����  $ %          � l ? 3       �  �  `�       Z       ��Q       ���� � ������������         ����  & '          � p B 6       �  &  �       Z       ��Q       ���� � ������������         ����  ) *          � t E 9       �  �  h�    
   Z       ��Q       ���� � ������������         ����  + ,          � x H <       �  R  �    	   Z	       ��Q       ���� � ������������          ����             � c 4 (       %  �  ��       [        ��R        ���� � ������������         ����             � h 7 +       2  ^  ��       [       ��R        ���� � ������������         ����    !          � m : .       >     ~�       [       ��R        ���� � ������������         ����  # $          � r = 1       K  �   j�       [       ��R       ���� � ������������         ����  % &          � w @ 4       W  z!  V�       [       ��R       ���� � ������������         ����  ' (          � | C 7       d  ."  B�       [       ��R       ���� � ������������         ����  ) *          � � F :       q  �"  .�       [       ��R       ���� � ������������         ����  + ,          � � I =       }  �#  �    	   [       ��R       ���� � ������������         ����  . /          � � L @       �  J$  �       [       ��R       ���� � ������������         ����  0 1          � � O C       �  �$  �      [	       ��R       ���� � ������������         ����  ! "          � { : .       /  �'  p>      \        ��S        ���� � �����  �           ����  # $          � � > 2       @  �(   E      \       ��S        ���� � �����  �           ����  % &          � � B 6       P  r)  �K      \       ��S        ���� � �����  �           ����  ( )          � � F :       a  D*   R      \       ��S       ���� � �����  �           ����  * +          � � J >       r  +  �X      \       ��S       ���� � �����  �           ����  , -          � � N B       �  �+  @_   	   \       ��S       ���� � �����  �           ����  . /          � � R F       �  �,  �e      \       ��S       ���� � �����  �           ����  0 1          � � V J       �  �-  `l      \       ��S       ���� � �����  �           ����  3 4          � � Z N       �  ^.  �r      \       ��S       ���� � �����  �           ����  5 6          � ^ R       �  0/  �y      \	       ��S       ���� � �����  �           ����  & '          � � J >       �  x2  8�      ]        ��T        ���� � �����  �            ����  ( )          � � N B       �  h3  ��      ]       ��T        ���� � �����  �            ����  * +          � � R F       �  X4  �      ]       ��T        ���� � �����  �            ����  - .          � V J       �  H5  ��   	   ]       ��T       ���� � �����  �            ����  / 0          � Z N       �  86  ��      ]       ��T       ���� � �����  �            ����  1 2          � ^ R       �  (7  h�      ]       ��T       ���� � �����  �            ����  3 4          � b V         8  ��      ]       ��T       ���� � �����  �            ����  5 6           � f Z       "  9  H      ]       ��T       ���� � �����  �            ����  8 9          '� j ^       7  �9  �	      ]       ��T       ���� � �����  �            ����  : ;          .� n b       M  �:  (      ]	       ��T       ���� � -  �  �            ����  + ,          � Y M       D  �>  �r      ^      	  ��U        ����	 � �����  �  !         ����  - .          � ] Q       _  �?  }   
   ^     	  ��U        ����	 � �����  �  !         ����  / 0          &� a U       z  �@  ��      ^     	  ��U        ����	 � �����  �  !         ����  2 3          -� e Y       �  �A  4�      ^     	  ��U       ����	 � �����  �  !         ����  4 5          4� i ]       �  �B  ��      ^     	  ��U       ����	 � �����  �  !         ����  6 7          ;� m a       �  �C  L�      ^     	  ��U       ����	 � �����  �  !         ����  8 9          B� q e       �  �D  ر      ^     	  ��U       ����	 � �����  �  !         ����  : ;          I� u i         
F  d�      ^     	  ��U       ����	 � �����  �  !         ����  = >          P� y m         G  ��       ^     	  ��U       ����	 � �����  �  !         ����  ? @          W� } q       7  &H  |�   ��  ^	     	  ��U       ����	 � 7  �  �  !          ����             ' D � '       b    H�       k        ��V        ���� � ������������"         ����             * H � *       k  �  ̍       k       ��V        ���� � ������������"         ����             - L � -       t  8  P�       k       ��V        ���� � ������������"         ����             0 P � 0       }  �  Ԕ       k       ��V       ���� � ������������"         ����             3 T � 3       �  d  X�       k       ��V       ���� � ������������"         ����             6 X � 6       �  �  ܛ       k       ��V       ���� � ������������"         ����              9 \ � 9       �  �  `�       k       ��V       ���� � ������������"         ����  ! "          < ` � <       �  &  �       k       ��V       ���� � ������������"         ����  # $          ? d � ?       �  �  h�    
   k       ��V       ���� � ������������"         ����  % &          B h � B       �  R  �    	   k	       ��V       ���� � ������������"          ����             . S � .       %  �  ��       l        ��W        ���� � ������������#         ����             2 W � 1       2  ^  ��       l       ��W        ���� � ������������#         ����             6 [ � 4       >     ~�       l       ��W        ���� � ������������#         ����             : _ � 7       K  �   j�       l       ��W       ���� � ������������#         ����             > c � :       W  z!  V�       l       ��W       ���� � ������������#         ����  ! "          B g � =       d  ."  B�       l       ��W       ���� � ������������#         ����  # $          F k � @       q  �"  .�       l       ��W       ���� � ������������#         ����  % &          J o � C       }  �#  �    	   l       ��W       ���� � ������������#         ����  ' (          N s � F       �  J$  �       l       ��W       ���� � ������������#         ����  ) *          R w � I       �  �$  �      l	       ��W       ���� � ������������#         ����             > b � 4       /  �'  p>      m        ��X        ���� � �����  �  $         ����             B g � 8       @  �(   E      m       ��X        ���� � �����  �  $         ����             F l � <       P  r)  �K      m       ��X        ���� � �����  �  $         ����    !          J q � @       a  D*   R      m       ��X       ���� � �����  �  $         ����  " #          N v � D       r  +  �X      m       ��X       ���� � �����  �  $         ����  $ %          R { � H       �  �+  @_   	   m       ��X       ���� � �����  �  $         ����  ' (          V � � L       �  �,  �e      m       ��X       ���� � �����  �  $         ����  ) *          Z � � P       �  �-  `l      m       ��X       ���� � �����  �  $         ����  + ,          ^ � � T       �  ^.  �r      m       ��X       ���� � �����  �  $         ����  - .          b � � X       �  0/  �y      m	       ��X       ���� � �����  �  $         ����             N z � D       �  x2  8�      n        ��Y        ���� � �����  �  %         ����    !          R  � H       �  h3  ��      n       ��Y        ���� � �����  �  %         ����  " #          V � � L       �  X4  �      n       ��Y        ���� � �����  �  %         ����  $ %          Z � � P       �  H5  ��   	   n       ��Y       ���� � �����  �  %         ����  & '          ^ � T       �  86  ��      n       ��Y       ���� � �����  �  %         ����  ( )          b � X       �  (7  h�      n       ��Y       ���� � �����  �  %         ����  + ,          f � \         8  ��      n       ��Y       ���� � �����  �  %         ����  - .          j � `       "  9  H      n       ��Y       ���� � �����  �  %         ����  / 0          n �  d       7  �9  �	      n       ��Y       ���� � �����  �  %         ����  1 2          r � 'h       M  �:  (      n	       ��Y       ���� � -  �  �  %         ����  " #          ] � S       D  �>  �r      o      	  ��Z        ����	 � �����  �  &         ����  $ %          a � W       _  �?  }   
   o     	  ��Z        ����	 � �����  �  &         ����  & '          e � [       z  �@  ��      o     	  ��Z        ����	 � �����  �  &         ����  ( )          i � &_       �  �A  4�      o     	  ��Z       ����	 � �����  �  &         ����  * +          m � -c       �  �B  ��      o     	  ��Z       ����	 � �����  �  &         ����  , -          q � 4g       �  �C  L�      o     	  ��Z       ����	 � �����  �  &         ����  / 0          u � ;k       �  �D  ر      o     	  ��Z       ����	 � �����  �  &         ����  1 2          y � Bo         
F  d�      o     	  ��Z       ����	 � �����  �  &         ����  3 4          } � Is         G  ��       o     	  ��Z       ����	 � �����  �  &         ����  5 6          � � Pw       7  &H  |�   ��  o	     	  ��Z       ����	 � 7  �  �  &          ����                         !   �  /       x        ��[        ���� � ������������'          ����                         (   �  �       x       ��[        ���� � ������������'          ����                         )            x       ��[        ���� � ������������'          ����                           )   *  T       x       ��[       ���� � ������������'          ����  	 
          $   $         *   H  �       x       ��[       ���� � ������������'          ����             (   (         +   f  �       x       ��[       ���� � ������������'          ����             ,   ,         +   �         x       ��[       ���� � ������������'          ����             0   0         ,   �  D       x       ��[       ���� � ������������'          ����             4   4         ,   �  �       x       ��[       ���� � ������������'          ����             8   8         -   �  �       x	       ��[       ���� � ������������'          ����             &  &         G   V	         y        ��\        ���� � ������������(          ����             *  *         I   �	  �       y       ��\        ���� � ������������(          ����  	 
          .  .         K   �	  j       y       ��\        ���� � ������������(          ����             2  2         M   

         y       ��\       ���� � ������������(          ����             6  6         N   F
  �       y       ��\       ���� � ������������(          ����             :  :         P   �
  �       y       ��\       ���� � ������������(          ����             >  >         R   �
  :        y       ��\       ���� � ������������(          ����             B ! B         T   �
  �        y       ��\       ���� � ������������(          ����             F # F         V   6  �!       y       ��\       ���� � ������������(          ����             J % J         W   r  V"       y	       ��\       ���� � ������������(          ����  	 
          7  7        ~   b  �1       z        ��]        ���� � ������������)         ����             <  <        �   �  �2       z       ��]        ���� � ������������)         ����             A  A        �     X4       z       ��]        ���� � ������������)         ����             F  F        �   p  �5       z       ��]       ���� � ������������)         ����             K  K        �   �  (7       z       ��]       ���� � ������������)         ����             P   P "       �   $  �8       z       ��]       ���� � ������������)         ����             U # U %       �   ~  �9       z       ��]       ���� � ������������)         ����             Z & Z (       �   �  `;       z       ��]       ���� � ������������)         ����             _ ) _ +       �   2  �<       z       ��]       ���� � ������������)         ����             d , d .       �   �  0>       z	       ��]       ���� � ������������)          ����             Q  Q        �   �  �T       {        ��^        ���� � ������������*         ����             V  V        �   l  W       {       ��^        ���� � ������������*         ����             [  [ !       �   �  tY       {       ��^        ���� � ������������*         ����             ` " ` $       �   \  �[       {       ��^       ���� � ������������*         ����             e % e '       �   �  $^       {       ��^       ���� � ������������*         ����             j ( j *       �   L  |`       {       ��^       ���� � ������������*         ����             o + o -       �   �  �b       {       ��^       ���� � ������������*         ����             t . t 0         <  ,e       {       ��^       ���� � ������������*         ����             y 1 y 3       	  �  �g       {       ��^       ���� � ������������*         ����    !          ~ 4 ~ 6         ,  �i       {	       ��^       ���� � ������������*          ����             j   j "       b    H�       |        ��_        ���� � ������������+         ����             o # o %       k  �  ̍       |       ��_        ���� � ������������+         ����             t & t (       t  8  P�       |       ��_        ���� � ������������+         ����             y ) y +       }  �  Ԕ       |       ��_       ���� � ������������+         ����             ~ , ~ .       �  d  X�       |       ��_       ���� � ������������+         ����             � / � 1       �  �  ܛ       |       ��_       ���� � ������������+         ����             � 2 � 4       �  �  `�       |       ��_       ���� � ������������+         ����    !          � 5 � 7       �  &  �       |       ��_       ���� � ������������+         ����  " #          � 8 � :       �  �  h�    
   |       ��_       ���� � ������������+         ����  $ %          � ; � =       �  R  �    	   |	       ��_       ���� � ������������+          ����             � ' � )       %  �  ��       }        ��`        ���� � ������������,         ����             � * � ,       2  ^  ��       }       ��`        ���� � ������������,         ����             � - � /       >     ~�       }       ��`        ���� � ������������,         ����             � 0 � 2       K  �   j�       }       ��`       ���� � ������������,         ����             � 3 � 5       W  z!  V�       }       ��`       ���� � ������������,         ����    !          � 6 � 8       d  ."  B�       }       ��`       ���� � ������������,         ����  " #          � 9 � ;       q  �"  .�       }       ��`       ���� � ������������,         ����  $ %          � < � >       }  �#  �    	   }       ��`       ���� � ������������,         ����  & '          � ? � A       �  J$  �       }       ��`       ���� � ������������,         ����  ( )          � B � D       �  �$  �      }	       ��`       ���� � ������������,         ����             � - � /       /  �'  p>      ~        ��a        ���� � �����  �  -         ����             � 1 � 3       @  �(   E      ~       ��a        ���� � �����  �  -         ����             � 5 � 7       P  r)  �K      ~       ��a        ���� � �����  �  -         ����              � 9 � ;       a  D*   R      ~       ��a       ���� � �����  �  -         ����  ! "          � = � ?       r  +  �X      ~       ��a       ���� � �����  �  -         ����  $ %          � A � C       �  �+  @_   	   ~       ��a       ���� � �����  �  -         ����  & '          � E � G       �  �,  �e      ~       ��a       ���� � �����  �  -         ����  ( )          � I � K       �  �-  `l      ~       ��a       ���� � �����  �  -         ����  * +          � M � O       �  ^.  �r      ~       ��a       ���� � �����  �  -         ����  , -          � Q � S       �  0/  �y      ~	       ��a       ���� � �����  �  -         ����             � = � ?       �  x2  8�              ��b        ���� � �����  �  .         ����              � A � C       �  h3  ��             ��b        ���� � �����  �  .         ����  ! "          � E � G       �  X4  �             ��b        ���� � �����  �  .         ����  # $          � I � K       �  H5  ��   	          ��b       ���� � �����  �  .         ����  % &          � M � O       �  86  ��             ��b       ���� � �����  �  .         ����  ' (          � Q � S       �  (7  h�             ��b       ���� � �����  �  .         ����  * +          � U � W         8  ��             ��b       ���� � �����  �  .         ����  , -          � Y � [       "  9  H             ��b       ���� � �����  �  .         ����  . /          � ] � _       7  �9  �	             ��b       ���� � �����  �  .         ����  0 1          � a � c       M  �:  (      	       ��b       ���� � -  �  �  .         ����  ! "          � L � N       D  �>  �r      �      	  ��c        ����	 � �����  �  /         ����  # $          � P � R       _  �?  }   
   �     	  ��c        ����	 � �����  �  /         ����  % &          � T � V       z  �@  ��      �     	  ��c        ����	 � �����  �  /         ����  ' (          � X � Z       �  �A  4�      �     	  ��c       ����	 � �����  �  /         ����  ) *          � \ � ^       �  �B  ��      �     	  ��c       ����	 � �����  �  /         ����  + ,          � ` � b       �  �C  L�      �     	  ��c       ����	 � �����  �  /         ����  . /           d  f       �  �D  ر      �     	  ��c       ����	 � �����  �  /         ����  0 1          h j         
F  d�      �     	  ��c       ����	 � �����  �  /         ����  2 3          l n         G  ��       �     	  ��c       ����	 � �����  �  /         ����  4 5          p r       7  &H  |�   ��  �	     	  ��c       ����	 � 7  �  �  /         ����             � T - !       J  |  �       �        ��d        ���� � ������������0         ����             � X 0 $       S    l�       �       ��d        ���� � ������������0         ����             � \ 3 '       \  �  ��       �       ��d        ���� � ������������0         ����  ! "          � ` 6 *       e  >  t�       �       ��d       ���� � ������������0         ����  # $          � d 9 -       n  �  ��       �       ��d       ���� � ������������0         ����  % &          � h < 0       w  j  |�       �       ��d       ���� � ������������0         ����  ' (          � l ? 3       �      �       �       ��d       ���� � ������������0         ����  ) *          � p B 6       �  �  ��       �       ��d       ���� � ������������0         ����  , -          � t E 9       �  ,  �    
   �       ��d       ���� � ������������0         ����  . /          � x H <       �  �  ��    	   �	       ��d       ���� � ������������0         ����              � c 4 (       	    ��       �        ��e        ���� � ������������1         ����  ! "          � h 7 +         �  ��       �       ��e        ���� � ������������1         ����  # $          � m : .       "  �  ��       �       ��e        ���� � ������������1         ����  & '          � r = 1       /  6  z�       �       ��e       ���� � ������������1         ����  ( )          � w @ 4       ;  �  f�       �       ��e       ���� � ������������1         ����  * +          � | C 7       H  �   R�       �       ��e       ���� � ������������1         ����  , -          � � F :       U  R!  >�       �       ��e       ���� � ������������1         ����  . /          � � I =       a  "  *�    	   �       ��e       ���� � ������������1         ����  1 2          � L @       n  �"  �       �       ��e       ���� � ������������1         ����  3 4          � O C       z  n#  �       �	       ��e       ���� � ������������1         ����  $ %          � { : .         >&  �1      �        ��f        ���� � �����  �  2         ����  & '          � � > 2          '  �8      �       ��f        ���� � �����  �  2         ����  ( )          � B 6       0  �'  ?      �       ��f        ���� � �����  �  2         ����  + ,          � F :       A  �(  �E      �       ��f       ���� � �����  �  2         ����  - .          � J >       R  �)  0L      �       ��f       ���� � �����  �  2         ����  / 0          � N B       c  X*  �R   	   �       ��f       ���� � �����  �  2         ����  1 2          � R F       t  *+  PY      �       ��f       ���� � �����  �  2         ����  3 4           � V J       �  �+  �_      �       ��f       ���� � �����  �  2         ����  6 7          &� Z N       �  �,  pf      �       ��f       ���� � �����  �  2         ����  8 9          ,� ^ R       �  �-   m      �	       ��f       ���� � �����  �  2         ����  ) *          � J >       f  �0  (�      �        ��g        ���� � �����  �  3         ����  + ,          � N B       |  �1  ��      �       ��g        ���� � �����  �  3         ����  - .          $� R F       �  �2  �      �       ��g        ���� � �����  �  3         ����  0 1          +� V J       �  �3  x�   	   �       ��g       ���� � �����  �  3         ����  2 3          2� Z N       �  �4  ��      �       ��g       ���� � �����  �  3         ����  4 5          9� ^ R       �  �5  X�      �       ��g       ���� � �����  �  3         ����  6 7          @� b V       �  �6  ��      �       ��g       ���� � �����  �  3         ����  8 9          G� f Z       �  x7  8�      �       ��g       ���� � �����  �  3         ����  ; <          N� j ^         h8  ��      �       ��g       ���� � �����  �  3         ����  = >          U� n b       )  X9        �	       ��g       ���� � -  �  �  3         ����  . /          ?� Y M         =  �b      �        ��h        ����	 � �����  �  4         ����  0 1          F� ] Q       7  &>  |m   
   �       ��h        ����	 � �����  �  4         ����  2 3          M� a U       R  4?  x      �       ��h        ����	 � �����  �  4         ����  5 6          T� e Y       m  B@  ��      �       ��h       ����	 � �����  �  4         ����  7 8          [� i ]       �  PA   �      �       ��h       ����	 � �����  �  4         ����  9 :          b� m a       �  ^B  ��      �       ��h       ����	 � �����  �  4         ����  ; <          i� q e       �  lC  8�      �       ��h       ����	 � �����  �  4         ����  = >          p� u i       �  zD  Ĭ      �       ��h       ����	 � �����  �  4         ����  @ A          w� y m       �  �E  P�       �       ��h       ����	 � �����  �  4         ����  B C          ~� } q         �F  ��   ��  �	       ��h       ����	 � 7  �  �  4         ����             M k � '       J  |  �       �        ��i        ���� � ������������5         ����             P o � *       S    l�       �       ��i        ���� � ������������5         ����             S s � -       \  �  ��       �       ��i        ���� � ������������5         ����             V w � 0       e  >  t�       �       ��i       ���� � ������������5         ����             Y { � 3       n  �  ��       �       ��i       ���� � ������������5         ����             \  � 6       w  j  |�       �       ��i       ���� � ������������5         ����    !          _ � � 9       �      �       �       ��i       ���� � ������������5         ����  " #          b � � <       �  �  ��       �       ��i       ���� � ������������5         ����  $ %          e � � ?       �  ,  �    
   �       ��i       ���� � ������������5         ����  & '          h � � B       �  �  ��    	   �	       ��i       ���� � ������������5         ����             T z � .       	    ��       �        ��j        ���� � ������������6         ����             X ~ � 1         �  ��       �       ��j        ���� � ������������6         ����             \ � � 4       "  �  ��       �       ��j        ���� � ������������6         ����             ` � � 7       /  6  z�       �       ��j       ���� � ������������6         ����              d � � :       ;  �  f�       �       ��j       ���� � ������������6         ����  " #          h � � =       H  �   R�       �       ��j       ���� � ������������6         ����  $ %          l � � @       U  R!  >�       �       ��j       ���� � ������������6         ����  & '          p � � C       a  "  *�    	   �       ��j       ���� � ������������6         ����  ( )          t � � F       n  �"  �       �       ��j       ���� � ������������6         ����  * +          x � I       z  n#  �       �	       ��j       ���� � ������������6         ����             d � � 4         >&  �1      �        ��k        ���� � �����  �  7         ����             h � � 8          '  �8      �       ��k        ���� � �����  �  7         ����              l � � <       0  �'  ?      �       ��k        ���� � �����  �  7         ����  ! "          p � @       A  �(  �E      �       ��k       ���� � �����  �  7         ����  # $          t � D       R  �)  0L      �       ��k       ���� � �����  �  7         ����  % &          x � H       c  X*  �R   	   �       ��k       ���� � �����  �  7         ����  ( )          | � L       t  *+  PY      �       ��k       ���� � �����  �  7         ����  * +          � � P       �  �+  �_      �       ��k       ���� � �����  �  7         ����  , -          � � T       �  �,  pf      �       ��k       ���� � �����  �  7         ����  . /          � � %X       �  �-   m      �	       ��k       ���� � �����  �  7         ����              t � D       f  �0  (�      �        ��l        ���� � �����  �  8         ����  ! "          x � H       |  �1  ��      �       ��l        ���� � �����  �  8         ����  # $          | � L       �  �2  �      �       ��l        ���� � �����  �  8         ����  % &          � � $P       �  �3  x�   	   �       ��l       ���� � �����  �  8         ����  ' (          � � +T       �  �4  ��      �       ��l       ���� � �����  �  8         ����  ) *          � � 2X       �  �5  X�      �       ��l       ���� � �����  �  8         ����  , -          � � 9\       �  �6  ��      �       ��l       ���� � �����  �  8         ����  . /          � � @`       �  x7  8�      �       ��l       ���� � �����  �  8         ����  0 1          � � Gd         h8  ��      �       ��l       ���� � �����  �  8         ����  2 3          � � Nh       )  X9        �	       ��l       ���� � -  �  �  8         ����  # $          � � 8S         =  �b      �        ��m        ����	 � �����  �  9         ����  % &          � � ?W       7  &>  |m   
   �       ��m        ����	 � �����  �  9         ����  ' (          � � F[       R  4?  x      �       ��m        ����	 � �����  �  9         ����  ) *          � � M_       m  B@  ��      �       ��m       ����	 � �����  �  9         ����  + ,          � � Tc       �  PA   �      �       ��m       ����	 � �����  �  9         ����  - .          � � [g       �  ^B  ��      �       ��m       ����	 � �����  �  9         ����  0 1          � � bk       �  lC  8�      �       ��m       ����	 � �����  �  9         ����  2 3          � � io       �  zD  Ĭ      �       ��m       ����	 � �����  �  9         ����  4 5          � � ps       �  �E  P�       �       ��m       ����	 � �����  �  9         ����  6 7          � � ww         �F  ��   ��  �	       ��m       ����	 � 7  �  �  9          ����             ;   ;            @  �       �         ��n        ���� � ������������:          ����             ?   ?             ^  �       �        ��n        ���� � ������������:          ����             C   C         !   |  �       �        ��n        ���� � ������������:          ����   	          G   G         !   �  4       �        ��n       ���� � ������������:          ����  
           K   K         "   �  p       �        ��n       ���� � ������������:          ����             O   O         #   �  �       �        ��n       ���� � ������������:          ����             S   S         #   �  �       �        ��n       ���� � ������������:          ����             W   W         $     $       �        ��n       ���� � ������������:          ����             [   [         $   0  `       �        ��n       ���� � ������������:          ����             _   _         %   N  �       �	        ��n       ���� � ������������:          ����             M  M         ;   �  R       �        ��o        ���� � ������������;          ����   	          Q  Q         =            �       ��o        ���� � ������������;          ����  
           U  U         ?   >  �       �       ��o        ���� � ������������;          ����             Y  Y         A   z  n       �       ��o       ���� � ������������;          ����             ]  ]         B   �  "       �       ��o       ���� � ������������;          ����             a  a         D   �  �       �       ��o       ���� � ������������;          ����             e  e         F   .	  �       �       ��o       ���� � ������������;          ����             i ! i         H   j	  >       �       ��o       ���� � ������������;          ����             m # m         J   �	  �       �       ��o       ���� � ������������;          ����             q % q         K   �	  �       �	       ��o       ���� � ������������;         ����  
           ^  ^        n   �
  H+       �        ��p        ���� � ������������<         ����             c  c        r   ,  �,       �       ��p        ���� � ������������<         ����             h  h        v   �  .       �       ��p        ���� � ������������<         ����             m  m        y   �  �/       �       ��p       ���� � ������������<         ����             r  r        }   :  �0       �       ��p       ���� � ������������<         ����             w   w "       �   �  P2       �       ��p       ���� � ������������<         ����             | # | %       �   �  �3       �       ��p       ���� � ������������<         ����             � & � (       �   H   5       �       ��p       ���� � ������������<         ����             � ) � +       �   �  �6       �       ��p       ���� � ������������<         ����             � , � .       �   �  �7       �	       ��p       ���� � ������������<         ����             x  x        �   d  �L       �        ��q        ���� � ������������=         ����             }  }        �   �  LO       �       ��q        ���� � ������������=         ����             �  � !       �   T  �Q       �       ��q        ���� � ������������=         ����             � " � $       �   �  �S       �       ��q       ���� � ������������=         ����             � % � '       �   D  TV       �       ��q       ���� � ������������=         ����             � ( � *       �   �  �X       �       ��q       ���� � ������������=         ����             � + � -       �   4  [       �       ��q       ���� � ������������=         ����             � . � 0       �   �  \]       �       ��q       ���� � ������������=         ����              � 1 � 3       �   $  �_       �       ��q       ���� � ������������=         ����  ! "          � 4 � 6       �   �  b       �	       ��q       ���� � ������������=         ����             �   � "       J  |  �       �        ��r        ���� � ������������>         ����             � # � %       S    l�       �       ��r        ���� � ������������>         ����             � & � (       \  �  ��       �       ��r        ���� � ������������>         ����             � ) � +       e  >  t�       �       ��r       ���� � ������������>         ����             � , � .       n  �  ��       �       ��r       ���� � ������������>         ����             � / � 1       w  j  |�       �       ��r       ���� � ������������>         ����              � 2 � 4       �      �       �       ��r       ���� � ������������>         ����  ! "          � 5 � 7       �  �  ��       �       ��r       ���� � ������������>         ����  # $          � 8 � :       �  ,  �    
   �       ��r       ���� � ������������>         ����  % &          � ; � =       �  �  ��    	   �	       ��r       ���� � ������������>         ����             � ' � )       	    ��       �        ��s        ���� � ������������?         ����             � * � ,         �  ��       �       ��s        ���� � ������������?         ����             � - � /       "  �  ��       �       ��s        ���� � ������������?         ����             � 0 � 2       /  6  z�       �       ��s       ���� � ������������?         ����             � 3 � 5       ;  �  f�       �       ��s       ���� � ������������?         ����  ! "          � 6 � 8       H  �   R�       �       ��s       ���� � ������������?         ����  # $          � 9 � ;       U  R!  >�       �       ��s       ���� � ������������?         ����  % &          � < � >       a  "  *�    	   �       ��s       ���� � ������������?         ����  ' (          � ? � A       n  �"  �       �       ��s       ���� � ������������?         ����  ) *          � B � D       z  n#  �       �	       ��s       ���� � ������������?         ����             � - � /         >&  �1      �        ��t        ���� � �����  �  @         ����             � 1 � 3          '  �8      �       ��t        ���� � �����  �  @         ����             � 5 � 7       0  �'  ?      �       ��t        ���� � �����  �  @         ����    !          � 9 � ;       A  �(  �E      �       ��t       ���� � �����  �  @         ����  " #          � = � ?       R  �)  0L      �       ��t       ���� � �����  �  @         ����  $ %          � A � C       c  X*  �R   	   �       ��t       ���� � �����  �  @         ����  ' (          � E � G       t  *+  PY      �       ��t       ���� � �����  �  @         ����  ) *          � I � K       �  �+  �_      �       ��t       ���� � �����  �  @         ����  + ,          � M � O       �  �,  pf      �       ��t       ���� � �����  �  @         ����  - .          � Q � S       �  �-   m      �	       ��t       ���� � �����  �  @         ����             � = � ?       f  �0  (�      �        ��u        ���� � �����  �  A         ����    !          � A � C       |  �1  ��      �       ��u        ���� � �����  �  A         ����  " #          � E � G       �  �2  �      �       ��u        ���� � �����  �  A         ����  $ %          � I � K       �  �3  x�   	   �       ��u       ���� � �����  �  A         ����  & '          � M � O       �  �4  ��      �       ��u       ���� � �����  �  A         ����  ( )          Q S       �  �5  X�      �       ��u       ���� � �����  �  A         ����  + ,          U W       �  �6  ��      �       ��u       ���� � �����  �  A         ����  - .          Y [       �  x7  8�      �       ��u       ���� � �����  �  A         ����  / 0          ] _         h8  ��      �       ��u       ���� � �����  �  A         ����  1 2          a c       )  X9        �	       ��u       ���� � -  �  �  A         ����  " #          L N         =  �b      �        ��v        ����	 � �����  �  B         ����  $ %          	P 	R       7  &>  |m   
   �       ��v        ����	 � �����  �  B         ����  & '          T V       R  4?  x      �       ��v        ����	 � �����  �  B         ����  ( )          X Z       m  B@  ��      �       ��v       ����	 � �����  �  B         ����  * +          \ ^       �  PA   �      �       ��v       ����	 � �����  �  B         ����  , -          !` !b       �  ^B  ��      �       ��v       ����	 � �����  �  B         ����  / 0          'd 'f       �  lC  8�      �       ��v       ����	 � �����  �  B         ����  1 2          -h -j       �  zD  Ĭ      �       ��v       ����	 � �����  �  B         ����  3 4          3l 3n       �  �E  P�       �       ��v       ����	 � �����  �  B         ����  5 6          9p 9r         �F  ��   ��  �	       ��v       ����	 � 7  �  �  B          ����             � T - !       2  �  �w       &        ��w        ���� � ������������C         ����             � X 0 $       ;  �  {       &       ��w        ���� � ������������C         ����             � \ 3 '       D    �~       &       ��w        ���� � ������������C         ����              � ` 6 *       M  �  �       &       ��w       ���� � ������������C         ����  ! "          � d 9 -       V  D  ��       &       ��w       ���� � ������������C         ����  # $          � h < 0       _  �  �       &       ��w       ���� � ������������C         ����  % &          � l ? 3       h  p  ��       &       ��w       ���� � ������������C         ����  ' (          � p B 6       q    $�       &       ��w       ���� � ������������C         ����  * +          � t E 9       z  �  ��    
   &       ��w       ���� � ������������C         ����  , -          � x H <       �  2  ,�    	   &	       ��w       ���� � ������������C          ����             � c 4 (       �  �  ��       '        ��x        ���� � ������������D         ����              � h 7 +       �  >  ��       '       ��x        ���� � ������������D         ����  ! "          � m : .         �  ��       '       ��x        ���� � ������������D         ����  $ %          � r = 1         �  ��       '       ��x       ���� � ������������D         ����  & '          � w @ 4         Z  v�       '       ��x       ���� � ������������D         ����  ( )          � | C 7       ,    b�       '       ��x       ���� � ������������D         ����  * +          � � F :       9  �  N�       '       ��x       ���� � ������������D         ����  , -          � � I =       E  v   :�    	   '       ��x       ���� � ������������D         ����  / 0          � � L @       R  *!  &�       '       ��x       ���� � ������������D         ����  1 2          � � O C       ^  �!  �       '	       ��x       ���� � ������������D         ����  " #          � { : .       �  �$  p%      (        ��y        ���� � �����  �  E         ����  $ %          � � > 2          �%   ,      (       ��y        ���� � �����  �  E         ����  & '          � � B 6         R&  �2      (       ��y        ���� � �����  �  E         ����  ) *          � � F :       !  $'   9      (       ��y       ���� � �����  �  E         ����  + ,          � � J >       2  �'  �?      (       ��y       ���� � �����  �  E         ����  - .          � � N B       C  �(  @F   	   (       ��y       ���� � �����  �  E         ����  / 0           � R F       T  �)  �L      (       ��y       ���� � �����  �  E         ����  1 2          � V J       d  l*  `S      (       ��y       ���� � �����  �  E         ����  4 5          � Z N       u  >+  �Y      (       ��y       ���� � �����  �  E         ����  6 7          � ^ R       �  ,  �`      (	       ��y       ���� � �����  �  E         ����  ' (          � � J >       B  X/  �      )        ��z        ���� � �����  �  F         ����  ) *          � N B       X  H0  ��      )       ��z        ���� � �����  �  F         ����  + ,          
� R F       n  81  ��      )       ��z        ���� � �����  �  F         ����  . /          � V J       �  (2  h�   	   )       ��z       ���� � �����  �  F         ����  0 1          � Z N       �  3  ��      )       ��z       ���� � �����  �  F         ����  2 3          � ^ R       �  4  H�      )       ��z       ���� � �����  �  F         ����  4 5          &� b V       �  �4  ��      )       ��z       ���� � �����  �  F         ����  6 7          -� f Z       �  �5  (�      )       ��z       ���� � �����  �  F         ����  9 :          4� j ^       �  �6  ��      )       ��z       ���� � �����  �  F         ����  ; <          ;� n b         �7  �      )	       ��z       ���� � -  �  �  F         ����  , -          %� Y M       �  �;  PS      *      	  ��{        ����	 � �����  �  G         ����  . /          ,� ] Q         �<  �]   
   *     	  ��{        ����	 � �����  �  G         ����  0 1          3� a U       *  �=  hh      *     	  ��{        ����	 � �����  �  G         ����  3 4          :� e Y       E  �>  �r      *     	  ��{       ����	 � �����  �  G         ����  5 6          A� i ]       `  �?  �}      *     	  ��{       ����	 � �����  �  G         ����  7 8          H� m a       {  �@  �      *     	  ��{       ����	 � �����  �  G         ����  9 :          O� q e       �  �A  ��      *     	  ��{       ����	 � �����  �  G         ����  ; <          V� u i       �  �B  $�      *     	  ��{       ����	 � �����  �  G         ����  > ?          ]� y m       �  �C  ��       *     	  ��{       ����	 � �����  �  G         ����  @ A          d� } q       �  E  <�   ��  *	     	  ��{       ����	 � 7  �  �  G          ����             4 Q � '       2  �  �w       7        ��|        ���� � ������������H         ����             7 U � *       ;  �  {       7       ��|        ���� � ������������H         ����             : Y � -       D    �~       7       ��|        ���� � ������������H         ����             = ] � 0       M  �  �       7       ��|       ���� � ������������H         ����             @ a � 3       V  D  ��       7       ��|       ���� � ������������H         ����             C e � 6       _  �  �       7       ��|       ���� � ������������H         ����              F i � 9       h  p  ��       7       ��|       ���� � ������������H         ����  ! "          I m � <       q    $�       7       ��|       ���� � ������������H         ����  # $          L q � ?       z  �  ��    
   7       ��|       ���� � ������������H         ����  % &          O u � B       �  2  ,�    	   7	       ��|       ���� � ������������H          ����             ; ` � .       �  �  ��       8        ��}        ���� � ������������I         ����             ? d � 1       �  >  ��       8       ��}        ���� � ������������I         ����             C h � 4         �  ��       8       ��}        ���� � ������������I         ����             G l � 7         �  ��       8       ��}       ���� � ������������I         ����             K p � :         Z  v�       8       ��}       ���� � ������������I         ����  ! "          O t � =       ,    b�       8       ��}       ���� � ������������I         ����  # $          S x � @       9  �  N�       8       ��}       ���� � ������������I         ����  % &          W | � C       E  v   :�    	   8       ��}       ���� � ������������I         ����  ' (          [ � � F       R  *!  &�       8       ��}       ���� � ������������I         ����  ) *          _ � � I       ^  �!  �       8	       ��}       ���� � ������������I         ����             K o � 4       �  �$  p%      9        ��~        ���� � �����  �  J         ����             O t � 8          �%   ,      9       ��~        ���� � �����  �  J         ����             S y � <         R&  �2      9       ��~        ���� � �����  �  J         ����    !          W ~ � @       !  $'   9      9       ��~       ���� � �����  �  J         ����  " #          [ � � D       2  �'  �?      9       ��~       ���� � �����  �  J         ����  $ %          _ � � H       C  �(  @F   	   9       ��~       ���� � �����  �  J         ����  ' (          c � � L       T  �)  �L      9       ��~       ���� � �����  �  J         ����  ) *          g � � P       d  l*  `S      9       ��~       ���� � �����  �  J         ����  + ,          k � T       u  >+  �Y      9       ��~       ���� � �����  �  J         ����  - .          o � X       �  ,  �`      9	       ��~       ���� � �����  �  J         ����             [ � � D       B  X/  �      :        ��        ���� � �����  �  K         ����    !          _ � � H       X  H0  ��      :       ��        ���� � �����  �  K         ����  " #          c � L       n  81  ��      :       ��        ���� � �����  �  K         ����  $ %          g � 
P       �  (2  h�   	   :       ��       ���� � �����  �  K         ����  & '          k � T       �  3  ��      :       ��       ���� � �����  �  K         ����  ( )          o � X       �  4  H�      :       ��       ���� � �����  �  K         ����  + ,          s � \       �  �4  ��      :       ��       ���� � �����  �  K         ����  - .          w � &`       �  �5  (�      :       ��       ���� � �����  �  K         ����  / 0          { � -d       �  �6  ��      :       ��       ���� � �����  �  K         ����  1 2           � 4h         �7  �      :	       ��       ���� � -  �  �  K         ����  " #          j � S       �  �;  PS      ;      	  ���        ����	 � �����  �  L         ����  $ %          n � %W         �<  �]   
   ;     	  ���        ����	 � �����  �  L         ����  & '          r � ,[       *  �=  hh      ;     	  ���        ����	 � �����  �  L         ����  ( )          v � 3_       E  �>  �r      ;     	  ���       ����	 � �����  �  L         ����  * +          z � :c       `  �?  �}      ;     	  ���       ����	 � �����  �  L         ����  , -          ~ � Ag       {  �@  �      ;     	  ���       ����	 � �����  �  L         ����  / 0          � � Hk       �  �A  ��      ;     	  ���       ����	 � �����  �  L         ����  1 2          � � Oo       �  �B  $�      ;     	  ���       ����	 � �����  �  L         ����  3 4          � � Vs       �  �C  ��       ;     	  ���       ����	 � �����  �  L         ����  5 6          � � ]w       �  E  <�   ��  ;	     	  ���       ����	 � 7  �  �  L          ����             !   !            �  F       D        ���        ���� � ������������M          ����             %   %            �  �	       D       ���        ���� � ������������M          ����             )   )            �  �	       D       ���        ���� � ������������M          ����             -   -            
  
       D       ���       ���� � ������������M          ����  	 
          1   1            (  P
       D       ���       ���� � ������������M          ����             5   5            F  �
       D       ���       ���� � ������������M          ����             9   9            d  �
       D       ���       ���� � ������������M          ����             =   =            �         D       ���       ���� � ������������M          ����             A   A            �  @       D       ���       ���� � ������������M          ����             E   E            �  |       D	       ���       ���� � ������������M          ����             3  3         /   6  �       E        ���        ���� � ������������N          ����             7  7         1   r  V       E       ���        ���� � ������������N          ����  	 
          ;  ;         3   �  
       E       ���        ���� � ������������N          ����             ?  ?         5   �  �       E       ���       ���� � ������������N          ����             C  C         6   &  r       E       ���       ���� � ������������N          ����             G  G         8   b  &       E       ���       ���� � ������������N          ����             K  K         :   �  �       E       ���       ���� � ������������N          ����             O ! O         <   �  �       E       ���       ���� � ������������N          ����             S # S         >     B       E       ���       ���� � ������������N          ����             W % W         ?   R  �       E	       ���       ���� � ������������N          ����  	 
          D  D        ^   B	  %       F        ���        ���� � ������������O         ����             I  I        b   �	  p&       F       ���        ���� � ������������O         ����             N  N        f   �	  �'       F       ���        ���� � ������������O         ����             S  S        i   P
  @)       F       ���       ���� � ������������O         ����             X  X        m   �
  �*       F       ���       ���� � ������������O         ����             ]   ] "       p     ,       F       ���       ���� � ������������O         ����             b # b %       t   ^  x-       F       ���       ���� � ������������O         ����             g & g (       x   �  �.       F       ���       ���� � ������������O         ����             l ) l +       {     H0       F       ���       ���� � ������������O         ����             q , q .          l  �1       F	       ���       ���� � ������������O          ����             ^  ^        �   �  $E       G        ���        ���� � ������������P         ����             c  c        �   L  |G       G       ���        ���� � ������������P         ����             h  h !       �   �  �I       G       ���        ���� � ������������P         ����             m " m $       �   <  ,L       G       ���       ���� � ������������P         ����             r % r '       �   �  �N       G       ���       ���� � ������������P         ����             w ( w *       �   ,  �P       G       ���       ���� � ������������P         ����             | + | -       �   �  4S       G       ���       ���� � ������������P         ����             � . � 0       �     �U       G       ���       ���� � ������������P         ����             � 1 � 3       �   �  �W       G       ���       ���� � ������������P         ����    !          � 4 � 6       �     <Z       G	       ���       ���� � ������������P          ����             w   w "       2  �  �w       H        ���        ���� � ������������Q         ����             | # | %       ;  �  {       H       ���        ���� � ������������Q         ����             � & � (       D    �~       H       ���        ���� � ������������Q         ����             � ) � +       M  �  �       H       ���       ���� � ������������Q         ����             � , � .       V  D  ��       H       ���       ���� � ������������Q         ����             � / � 1       _  �  �       H       ���       ���� � ������������Q         ����             � 2 � 4       h  p  ��       H       ���       ���� � ������������Q         ����    !          � 5 � 7       q    $�       H       ���       ���� � ������������Q         ����  " #          � 8 � :       z  �  ��    
   H       ���       ���� � ������������Q         ����  $ %          � ; � =       �  2  ,�    	   H	       ���       ���� � ������������Q          ����             � ' � )       �  �  ��       I        ���        ���� � ������������R         ����             � * � ,       �  >  ��       I       ���        ���� � ������������R         ����             � - � /         �  ��       I       ���        ���� � ������������R         ����             � 0 � 2         �  ��       I       ���       ���� � ������������R         ����             � 3 � 5         Z  v�       I       ���       ���� � ������������R         ����    !          � 6 � 8       ,    b�       I       ���       ���� � ������������R         ����  " #          � 9 � ;       9  �  N�       I       ���       ���� � ������������R         ����  $ %          � < � >       E  v   :�    	   I       ���       ���� � ������������R         ����  & '          � ? � A       R  *!  &�       I       ���       ���� � ������������R         ����  ( )          � B � D       ^  �!  �       I	       ���       ���� � ������������R         ����             � - � /       �  �$  p%      J        ���        ���� � �����  �  S         ����             � 1 � 3          �%   ,      J       ���        ���� � �����  �  S         ����             � 5 � 7         R&  �2      J       ���        ���� � �����  �  S         ����              � 9 � ;       !  $'   9      J       ���       ���� � �����  �  S         ����  ! "          � = � ?       2  �'  �?      J       ���       ���� � �����  �  S         ����  $ %          � A � C       C  �(  @F   	   J       ���       ���� � �����  �  S         ����  & '          � E � G       T  �)  �L      J       ���       ���� � �����  �  S         ����  ( )          � I � K       d  l*  `S      J       ���       ���� � �����  �  S         ����  * +          � M � O       u  >+  �Y      J       ���       ���� � �����  �  S         ����  , -          � Q � S       �  ,  �`      J	       ���       ���� � �����  �  S         ����             � = � ?       B  X/  �      K        ���        ���� � �����  �  T         ����              � A � C       X  H0  ��      K       ���        ���� � �����  �  T         ����  ! "          � E � G       n  81  ��      K       ���        ���� � �����  �  T         ����  # $          � I � K       �  (2  h�   	   K       ���       ���� � �����  �  T         ����  % &          � M � O       �  3  ��      K       ���       ���� � �����  �  T         ����  ' (          � Q � S       �  4  H�      K       ���       ���� � �����  �  T         ����  * +          � U � W       �  �4  ��      K       ���       ���� � �����  �  T         ����  , -          � Y � [       �  �5  (�      K       ���       ���� � �����  �  T         ����  . /          � ] � _       �  �6  ��      K       ���       ���� � �����  �  T         ����  0 1          � a � c         �7  �      K	       ���       ���� � -  �  �  T         ����  ! "          � L � N       �  �;  PS      L      	  ���        ����	 � �����  �  U         ����  # $          � P � R         �<  �]   
   L     	  ���        ����	 � �����  �  U         ����  % &          � T � V       *  �=  hh      L     	  ���        ����	 � �����  �  U         ����  ' (          � X � Z       E  �>  �r      L     	  ���       ����	 � �����  �  U         ����  ) *          \ ^       `  �?  �}      L     	  ���       ����	 � �����  �  U         ����  + ,          ` b       {  �@  �      L     	  ���       ����	 � �����  �  U         ����  . /          d f       �  �A  ��      L     	  ���       ����	 � �����  �  U         ����  0 1          h j       �  �B  $�      L     	  ���       ����	 � �����  �  U         ����  2 3          l n       �  �C  ��       L     	  ���       ����	 � �����  �  U         ����  4 5          p r       �  E  <�   ��  L	     	  ���       ����	 � 7  �  �  U         ����             � T - !       z  �  ��       �      �   �        ���� � ������������V         ����             � X 0 $       �  2  ,�       �     �   �        ���� � ������������V         ����             � \ 3 '       �  �  ��       �     �   �        ���� � ������������V         ����    !          � ` 6 *       �  ^  4�       �     �   �       ���� � ������������V         ����  " #          � d 9 -       �  �  ��       �     �   �       ���� � ������������V         ����  $ %          � h < 0       �  �  <�       �     �   �       ���� � ������������V         ����  & '          � l ? 3       �     ��       �     �   �       ���� � ������������V         ����  ( )          � p B 6       �  �  D�       �     �   �       ���� � ������������V         ����  + ,          � t E 9       �  L  ȯ    
   �     �   �       ���� � ������������V         ����  - .          � x H <       �  �  L�    	   �	     �   �       ���� � ������������V         ����             � c 4 (       A  :   ��       �      �   �        ���� � ������������W         ����    !          � h 7 +       N  �   ��       �     �   �        ���� � ������������W         ����  " #          � m : .       Z  �!  n�       �     �   �        ���� � ������������W         ����  % &          � r = 1       g  V"  Z�       �     �   �       ���� � ������������W         ����  ' (          � w @ 4       s  
#  F�       �     �   �       ���� � ������������W         ����  ) *          � | C 7       �  �#  2�       �     �   �       ���� � ������������W         ����  + ,          � � F :       �  r$  �       �     �   �       ���� � ������������W         ����  - .          � � I =       �  &%  
   	   �     �   �       ���� � ������������W         ����  0 1          � � L @       �  �%  �      �     �   �       ���� � ������������W         ����  2 3          � O C       �  �&  �      �	     �   �       ���� � ������������W         ����  # $          � { : .       O  ^)  �J      �      �   �        ���� � �����  �  X         ����  % &          � � > 2       `  0*  �Q      �     �   �        ���� � �����  �  X         ����  ' (          � � B 6       p  +  X      �     �   �        ���� � �����  �  X         ����  * +           � F :       �  �+  �^      �     �   �       ���� � �����  �  X         ����  , -          � J >       �  �,  0e      �     �   �       ���� � �����  �  X         ����  . /          � N B       �  x-  �k   	   �     �   �       ���� � �����  �  X         ����  0 1          � R F       �  J.  Pr      �     �   �       ���� � �����  �  X         ����  2 3          � V J       �  /  �x      �     �   �       ���� � �����  �  X         ����  5 6          � Z N       �  �/  p      �     �   �       ���� � �����  �  X         ����  7 8          $� ^ R       �  �0   �      �	     �   �       ���� � �����  �  X         ����  ( )          � J >       �  4  H�      �      �   �        ���� � �����  �  Y         ����  * +          � N B       �  �4  ��      �     �   �        ���� � �����  �  Y         ����  , -          � R F       �  �5  (�      �     �   �        ���� � �����  �  Y         ����  / 0          #� V J       �  �6  ��   	   �     �   �       ���� � �����  �  Y         ����  1 2          *� Z N         �7  �      �     �   �       ���� � �����  �  Y         ����  3 4          1� ^ R         �8  x�      �     �   �       ���� � �����  �  Y         ����  5 6          8� b V       0  �9  �      �     �   �       ���� � �����  �  Y         ����  7 8          ?� f Z       F  �:  X      �     �   �       ���� � �����  �  Y         ����  : ;          F� j ^       [  �;  �      �     �   �       ���� � �����  �  Y         ����  < =          M� n b       q  x<  8       �	     �   �       ���� � -  �  �  Y         ����  - .          7� Y M       l  8@  0�      �      �   �        ����	 � �����  �  Z         ����  / 0          >� ] Q       �  FA  ��   
   �     �   �        ����	 � �����  �  Z         ����  1 2          E� a U       �  TB  H�      �     �   �        ����	 � �����  �  Z         ����  4 5          L� e Y       �  bC  ԡ      �     �   �       ����	 � �����  �  Z         ����  6 7          S� i ]       �  pD  `�      �     �   �       ����	 � �����  �  Z         ����  8 9          Z� m a       �  ~E  �      �     �   �       ����	 � �����  �  Z         ����  : ;          a� q e         �F  x�      �     �   �       ����	 � �����  �  Z         ����  < =          h� u i       )  �G  �      �     �   �       ����	 � �����  �  Z         ����  ? @          o� y m       D  �H  ��       �     �   �       ����	 � �����  �  Z         ����  A B          v� } q       _  �I  �   ��  �	     �   �       ����	 � 7  �  �  Z         ����             E c � '       z  �  ��       �      �   �        ���� � ������������[         ����             H g � *       �  2  ,�       �     �   �        ���� � ������������[         ����             K k � -       �  �  ��       �     �   �        ���� � ������������[         ����             N o � 0       �  ^  4�       �     �   �       ���� � ������������[         ����             Q s � 3       �  �  ��       �     �   �       ���� � ������������[         ����             T w � 6       �  �  <�       �     �   �       ���� � ������������[         ����    !          W { � 9       �     ��       �     �   �       ���� � ������������[         ����  " #          Z  � <       �  �  D�       �     �   �       ���� � ������������[         ����  $ %          ] � � ?       �  L  ȯ    
   �     �   �       ���� � ������������[         ����  & '          ` � � B       �  �  L�    	   �	     �   �       ���� � ������������[         ����             L r � .       A  :   ��       �      �   �        ���� � ������������\         ����             P v � 1       N  �   ��       �     �   �        ���� � ������������\         ����             T z � 4       Z  �!  n�       �     �   �        ���� � ������������\         ����             X ~ � 7       g  V"  Z�       �     �   �       ���� � ������������\         ����              \ � � :       s  
#  F�       �     �   �       ���� � ������������\         ����  " #          ` � � =       �  �#  2�       �     �   �       ���� � ������������\         ����  $ %          d � � @       �  r$  �       �     �   �       ���� � ������������\         ����  & '          h � � C       �  &%  
   	   �     �   �       ���� � ������������\         ����  ( )          l � � F       �  �%  �      �     �   �       ���� � ������������\         ����  * +          p � � I       �  �&  �      �	     �   �       ���� � ������������\         ����             \ � � 4       O  ^)  �J      �      �   �        ���� � �����  �  ]         ����             ` � � 8       `  0*  �Q      �     �   �        ���� � �����  �  ]         ����              d � � <       p  +  X      �     �   �        ���� � �����  �  ]         ����  ! "          h � � @       �  �+  �^      �     �   �       ���� � �����  �  ]         ����  # $          l � � D       �  �,  0e      �     �   �       ���� � �����  �  ]         ����  % &          p � H       �  x-  �k   	   �     �   �       ���� � �����  �  ]         ����  ( )          t � L       �  J.  Pr      �     �   �       ���� � �����  �  ]         ����  * +          x � P       �  /  �x      �     �   �       ���� � �����  �  ]         ����  , -          | � T       �  �/  p      �     �   �       ���� � �����  �  ]         ����  . /          � � X       �  �0   �      �	     �   �       ���� � �����  �  ]         ����              l � D       �  4  H�      �      �   �        ���� � �����  �  ^         ����  ! "          p � H       �  �4  ��      �     �   �        ���� � �����  �  ^         ����  # $          t � L       �  �5  (�      �     �   �        ���� � �����  �  ^         ����  % &          x � P       �  �6  ��   	   �     �   �       ���� � �����  �  ^         ����  ' (          | � #T         �7  �      �     �   �       ���� � �����  �  ^         ����  ) *          � � *X         �8  x�      �     �   �       ���� � �����  �  ^         ����  , -          � � 1\       0  �9  �      �     �   �       ���� � �����  �  ^         ����  . /          � � 8`       F  �:  X      �     �   �       ���� � �����  �  ^         ����  0 1          � � ?d       [  �;  �      �     �   �       ���� � �����  �  ^         ����  2 3          � � Fh       q  x<  8       �	     �   �       ���� � -  �  �  ^         ����  # $          { � 0S       l  8@  0�      �      �   �        ����	 � �����  �  _         ����  % &           � 7W       �  FA  ��   
   �     �   �        ����	 � �����  �  _         ����  ' (          � � >[       �  TB  H�      �     �   �        ����	 � �����  �  _         ����  ) *          � � E_       �  bC  ԡ      �     �   �       ����	 � �����  �  _         ����  + ,          � � Lc       �  pD  `�      �     �   �       ����	 � �����  �  _         ����  - .          � � Sg       �  ~E  �      �     �   �       ����	 � �����  �  _         ����  0 1          � � Zk         �F  x�      �     �   �       ����	 � �����  �  _         ����  2 3          � � ao       )  �G  �      �     �   �       ����	 � �����  �  _         ����  4 5          � � hs       D  �H  ��       �     �   �       ����	 � �����  �  _         ����  6 7          � � ow       _  �I  �   ��  �	     �   �       ����	 � 7  �  �  _          ����             3   3         2   `	  �       �      �   �        ���� � ������������`          ����             7   7         0   ~	  �       �     �   �        ���� � ������������`          ����             ;   ;         1   �	  8       �     �   �        ���� � ������������`          ����   	          ?   ?         1   �	  t       �     �   �       ���� � ������������`          ����  
           C   C         2   �	  �       �     �   �       ���� � ������������`          ����             G   G         3   �	  �       �     �   �       ���� � ������������`          ����             K   K         3   
  (       �     �   �       ���� � ������������`          ����             O   O         4   2
  d       �     �   �       ���� � ������������`          ����             S   S         4   P
  �       �     �   �       ���� � ������������`          ����             W   W         5   n
  �       �	     �   �       ���� � ������������`          ����             E  E         S   �
  �        �      �   �        ���� � ������������a          ����   	          I  I         U   "  f!       �     �   �        ���� � ������������a          ����  
           M  M         W   ^  "       �     �   �        ���� � ������������a          ����             Q  Q         Y   �  �"       �     �   �       ���� � ������������a          ����             U  U         Z   �  �#       �     �   �       ���� � ������������a          ����             Y  Y         \     6$       �     �   �       ���� � ������������a          ����             ]  ]         ^   N  �$       �     �   �       ���� � ������������a          ����             a ! a         `   �  �%       �     �   �       ���� � ������������a          ����             e # e         b   �  R&       �     �   �       ���� � ������������a          ����             i % i         c     '       �	     �   �       ���� � ������������a         ����  
           V  V        �   �  �7       �      �   �        ���� � ������������b         ����             [  [        �   L  09       �     �   �        ���� � ������������b         ����             `  `        �   �  �:       �     �   �        ���� � ������������b         ����             e  e        �       <       �     �   �       ���� � ������������b         ����             j  j        �   Z  h=       �     �   �       ���� � ������������b         ����             o   o "       �   �  �>       �     �   �       ���� � ������������b         ����             t # t %       �     8@       �     �   �       ���� � ������������b         ����             y & y (       �   h  �A       �     �   �       ���� � ������������b         ����             ~ ) ~ +       �   �  C       �     �   �       ���� � ������������b         ����             � , � .       �     pD       �	     �   �       ���� � ������������b         ����             p  p        �   �  �\       �      �   �        ���� � ������������c         ����             u  u        �   �  �^       �     �   �        ���� � ������������c         ����             z  z !       �   t  Da       �     �   �        ���� � ������������c         ����              "  $       �   �  �c       �     �   �       ���� � ������������c         ����             � % � '         d  �e       �     �   �       ���� � ������������c         ����             � ( � *         �  Lh       �     �   �       ���� � ������������c         ����             � + � -         T  �j       �     �   �       ���� � ������������c         ����             � . � 0         �  �l       �     �   �       ���� � ������������c         ����              � 1 � 3         D  To       �     �   �       ���� � ������������c         ����  ! "          � 4 � 6       #  �  �q       �	     �   �       ���� � ������������c         ����             �   � "       z  �  ��       �      �   �        ���� � ������������d         ����             � # � %       �  2  ,�       �     �   �        ���� � ������������d         ����             � & � (       �  �  ��       �     �   �        ���� � ������������d         ����             � ) � +       �  ^  4�       �     �   �       ���� � ������������d         ����             � , � .       �  �  ��       �     �   �       ���� � ������������d         ����             � / � 1       �  �  <�       �     �   �       ���� � ������������d         ����              � 2 � 4       �     ��       �     �   �       ���� � ������������d         ����  ! "          � 5 � 7       �  �  D�       �     �   �       ���� � ������������d         ����  # $          � 8 � :       �  L  ȯ    
   �     �   �       ���� � ������������d         ����  % &          � ; � =       �  �  L�    	   �	     �   �       ���� � ������������d         ����             � ' � )       A  :   ��       �      �   �        ���� � ������������e         ����             � * � ,       N  �   ��       �     �   �        ���� � ������������e         ����             � - � /       Z  �!  n�       �     �   �        ���� � ������������e         ����             � 0 � 2       g  V"  Z�       �     �   �       ���� � ������������e         ����             � 3 � 5       s  
#  F�       �     �   �       ���� � ������������e         ����  ! "          � 6 � 8       �  �#  2�       �     �   �       ���� � ������������e         ����  # $          � 9 � ;       �  r$  �       �     �   �       ���� � ������������e         ����  % &          � < � >       �  &%  
   	   �     �   �       ���� � ������������e         ����  ' (          � ? � A       �  �%  �      �     �   �       ���� � ������������e         ����  ) *          � B � D       �  �&  �      �	     �   �       ���� � ������������e         ����             � - � /       O  ^)  �J      �      �   �        ���� � �����  �  f         ����             � 1 � 3       `  0*  �Q      �     �   �        ���� � �����  �  f         ����             � 5 � 7       p  +  X      �     �   �        ���� � �����  �  f         ����    !          � 9 � ;       �  �+  �^      �     �   �       ���� � �����  �  f         ����  " #          � = � ?       �  �,  0e      �     �   �       ���� � �����  �  f         ����  $ %          � A � C       �  x-  �k   	   �     �   �       ���� � �����  �  f         ����  ' (          � E � G       �  J.  Pr      �     �   �       ���� � �����  �  f         ����  ) *          � I � K       �  /  �x      �     �   �       ���� � �����  �  f         ����  + ,          � M � O       �  �/  p      �     �   �       ���� � �����  �  f         ����  - .          � Q � S       �  �0   �      �	     �   �       ���� � �����  �  f         ����             � = � ?       �  4  H�      �      �   �        ���� � �����  �  g         ����    !          � A � C       �  �4  ��      �     �   �        ���� � �����  �  g         ����  " #          � E � G       �  �5  (�      �     �   �        ���� � �����  �  g         ����  $ %          � I � K       �  �6  ��   	   �     �   �       ���� � �����  �  g         ����  & '          � M � O         �7  �      �     �   �       ���� � �����  �  g         ����  ( )          � Q � S         �8  x�      �     �   �       ���� � �����  �  g         ����  + ,          � U � W       0  �9  �      �     �   �       ���� � �����  �  g         ����  - .          Y [       F  �:  X      �     �   �       ���� � �����  �  g         ����  / 0          ] _       [  �;  �      �     �   �       ���� � �����  �  g         ����  1 2          a c       q  x<  8       �	     �   �       ���� � -  �  �  g         ����  " #          � L � N       l  8@  0�      �      �   �        ����	 � �����  �  h         ����  $ %          P R       �  FA  ��   
   �     �   �        ����	 � �����  �  h         ����  & '          T V       �  TB  H�      �     �   �        ����	 � �����  �  h         ����  ( )          X Z       �  bC  ԡ      �     �   �       ����	 � �����  �  h         ����  * +          \ ^       �  pD  `�      �     �   �       ����	 � �����  �  h         ����  , -          ` b       �  ~E  �      �     �   �       ����	 � �����  �  h         ����  / 0          d f         �F  x�      �     �   �       ����	 � �����  �  h         ����  1 2          %h %j       )  �G  �      �     �   �       ����	 � �����  �  h         ����  3 4          +l +n       D  �H  ��       �     �   �       ����	 � �����  �  h         ����  5 6          1p 1r       _  �I  �   ��  �	     �   �       ����	 � 7  �  �  h         ����	              � T - !       ����L  ȯ       �      �� ���        ���� � ������������i         ����	              � X 0 $       �����  L�       �     �� ���        ���� � ������������i         ����	              � \ 3 '       ����x  ж       �     �� ���        ���� � ������������i         ����	              � ` 6 *       ����  T�       �     �� ���       ���� � ������������i         ����	    !           � d 9 -       �����  ؽ       �     �� ���       ���� � ������������i         ����	  " #           � h < 0       ����:   \�       �     �� ���       ���� � ������������i         ����	  $ %           � l ? 3       �����   ��       �     �� ���       ���� � ������������i         ����	  & '           � p B 6       ����f!  d�       �     �� ���       ���� � ������������i         ����	  ) *           � t E 9       �����!  ��    
   �     �� ���       ���� � ������������i         ����	  + ,           � x H <       �����"  l�    	   �	     �� ���       ���� � ������������i         ����	              � c 4 (       �����$  f      �      �� ���        ���� � ������������j         ����	              � h 7 +       �����%  R      �     �� ���        ���� � ������������j         ����	    !           � m : .       ����R&  >      �     �� ���        ���� � ������������j         ����	  # $           � r = 1       ����'  *      �     �� ���       ���� � ������������j         ����	  % &           � w @ 4       �����'        �     �� ���       ���� � ������������j         ����	  ' (           � | C 7       ����n(        �     �� ���       ���� � ������������j         ����	  ) *           � � F :       ����")  �      �     �� ���       ���� � ������������j         ����	  + ,           � � I =       �����)  �$   	   �     �� ���       ���� � ������������j         ����	  . /           � � L @       �����*  �)      �     �� ���       ���� � ������������j         ����	  0 1           � � O C       ����>+  �.      �	     �� ���       ���� � ������������j         ����	  ! "           � { : .       ����.  pp      �      �� ���        ���� � �����  �  k         ����	  # $           � � > 2       �����.   w      �     �� ���        ���� � �����  �  k         ����	  % &           � � B 6       �����/  �}      �     �� ���        ���� � �����  �  k         ����	  ( )           � � F :       �����0   �      �     �� ���       ���� � �����  �  k         ����	  * +           � � J >       ����V1  ��      �     �� ���       ���� � �����  �  k         ����	  , -           � � N B       ����(2  @�   	   �     �� ���       ���� � �����  �  k         ����	  . /           � � R F       �����2  З      �     �� ���       ���� � �����  �  k         ����	  0 1           � V J       �����3  `�      �     �� ���       ���� � �����  �  k         ����	  3 4           � Z N       �����4  �      �     �� ���       ���� � �����  �  k         ����	  5 6           � ^ R       ����p5  ��      �	     �� ���       ���� � �����  �  k         ����	  & '           � � J >       �����8  x�      �      �� ���        ���� � �����  �  l         ����	  ( )           � � N B       �����9  �      �     �� ���        ���� � �����  �  l         ����	  * +           � R F       �����:  X      �     �� ���        ���� � �����  �  l         ����	  - .           � V J       �����;  �   	   �     �� ���       ���� � �����  �  l         ����	  / 0           � Z N       ����x<  8       �     �� ���       ���� � �����  �  l         ����	  1 2           � ^ R       ����h=  �(      �     �� ���       ���� � �����  �  l         ����	  3 4           !� b V       ����X>  1      �     �� ���       ���� � �����  �  l         ����	  5 6           (� f Z       ����H?  �9      �     �� ���       ���� � �����  �  l         ����	  8 9           /� j ^       ����8@  �A      �     �� ���       ���� � �����  �  l         ����	  : ;           6� n b       ����(A  hJ      �	     �� ���       ���� � �����  �  l         ����	  + ,            � Y M       �����D  �      �      �� ���        ����	 � �����  �  m         ����	  - .           '� ] Q       �����E  ��   
   �     �� ���        ����	 � �����  �  m         ����	  / 0           .� a U       ����G  (�      �     �� ���        ����	 � �����  �  m         ����	  2 3           5� e Y       ����H  ��      �     �� ���       ����	 � �����  �  m         ����	  4 5           <� i ]       ���� I  @�      �     �� ���       ����	 � �����  �  m         ����	  6 7           C� m a       ����.J  ��      �     �� ���       ����	 � �����  �  m         ����	  8 9           J� q e       ����<K  X�      �     �� ���       ����	 � �����  �  m         ����	  : ;           Q� u i       ����JL  ��      �     �� ���       ����	 � �����  �  m         ����	  = >           X� y m       ����XM  p       �     �� ���       ����	 � �����  �  m         ����	  ? @           _� } q       ����fN  �   ��  �	     �� ���       ����	 � �����  �  m         ����	              / L � '       ����L  ȯ       �      �� ���        ���� � ������������n         ����	              2 P � *       �����  L�       �     �� ���        ���� � ������������n         ����	              5 T � -       ����x  ж       �     �� ���        ���� � ������������n         ����	              8 X � 0       ����  T�       �     �� ���       ���� � ������������n         ����	              ; \ � 3       �����  ؽ       �     �� ���       ���� � ������������n         ����	              > ` � 6       ����:   \�       �     �� ���       ���� � ������������n         ����	               A d � 9       �����   ��       �     �� ���       ���� � ������������n         ����	  ! "           D h � <       ����f!  d�       �     �� ���       ���� � ������������n         ����	  # $           G l � ?       �����!  ��    
   �     �� ���       ���� � ������������n         ����	  % &           J p � B       �����"  l�    	   �	     �� ���       ���� � ������������n         ����	              6 [ � .       �����$  f      �      �� ���        ���� � ������������o         ����	              : _ � 1       �����%  R      �     �� ���        ���� � ������������o         ����	              > c � 4       ����R&  >      �     �� ���        ���� � ������������o         ����	              B g � 7       ����'  *      �     �� ���       ���� � ������������o         ����	              F k � :       �����'        �     �� ���       ���� � ������������o         ����	  ! "           J o � =       ����n(        �     �� ���       ���� � ������������o         ����	  # $           N s � @       ����")  �      �     �� ���       ���� � ������������o         ����	  % &           R w � C       �����)  �$   	   �     �� ���       ���� � ������������o         ����	  ' (           V { � F       �����*  �)      �     �� ���       ���� � ������������o         ����	  ) *           Z  � I       ����>+  �.      �	     �� ���       ���� � ������������o         ����	              F j � 4       ����.  pp      �      �� ���        ���� � �����  �  p         ����	              J o � 8       �����.   w      �     �� ���        ���� � �����  �  p         ����	              N t � <       �����/  �}      �     �� ���        ���� � �����  �  p         ����	    !           R y � @       �����0   �      �     �� ���       ���� � �����  �  p         ����	  " #           V ~ � D       ����V1  ��      �     �� ���       ���� � �����  �  p         ����	  $ %           Z � � H       ����(2  @�   	   �     �� ���       ���� � �����  �  p         ����	  ' (           ^ � � L       �����2  З      �     �� ���       ���� � �����  �  p         ����	  ) *           b � � P       �����3  `�      �     �� ���       ���� � �����  �  p         ����	  + ,           f �  T       �����4  �      �     �� ���       ���� � �����  �  p         ����	  - .           j � X       ����p5  ��      �	     �� ���       ���� � �����  �  p         ����	              V � � D       �����8  x�      �      �� ���        ���� � �����  �  q         ����	    !           Z � � H       �����9  �      �     �� ���        ���� � �����  �  q         ����	  " #           ^ � � L       �����:  X      �     �� ���        ���� � �����  �  q         ����	  $ %           b � P       �����;  �   	   �     �� ���       ���� � �����  �  q         ����	  & '           f � T       ����x<  8       �     �� ���       ���� � �����  �  q         ����	  ( )           j � X       ����h=  �(      �     �� ���       ���� � �����  �  q         ����	  + ,           n � \       ����X>  1      �     �� ���       ���� � �����  �  q         ����	  - .           r � !`       ����H?  �9      �     �� ���       ���� � �����  �  q         ����	  / 0           v � (d       ����8@  �A      �     �� ���       ���� � �����  �  q         ����	  1 2           z � /h       ����(A  hJ      �	     �� ���       ���� � �����  �  q         ����	  " #           e � S       �����D  �      �      �� ���        ����	 � �����  �  r         ����	  $ %           i �  W       �����E  ��   
   �     �� ���        ����	 � �����  �  r         ����	  & '           m � '[       ����G  (�      �     �� ���        ����	 � �����  �  r         ����	  ( )           q � ._       ����H  ��      �     �� ���       ����	 � �����  �  r         ����	  * +           u � 5c       ���� I  @�      �     �� ���       ����	 � �����  �  r         ����	  , -           y � <g       ����.J  ��      �     �� ���       ����	 � �����  �  r         ����	  / 0           } � Ck       ����<K  X�      �     �� ���       ����	 � �����  �  r         ����	  1 2           � � Jo       ����JL  ��      �     �� ���       ����	 � �����  �  r         ����	  3 4           � � Qs       ����XM  p       �     �� ���       ����	 � �����  �  r         ����	  5 6           � � Xw       ����fN  �   ��  �	     �� ���       ����	 � �����  �  r          ����	                          ����  .J       �      �� ���        ���� � ������������s          ����	                            ����.  \       �     �� ���        ���� � ������������s          ����	              $   $         ����L  �       �     �� ���        ���� � ������������s          ����	              (   (         ����j  �       �     �� ���       ���� � ������������s          ����	  	 
           ,   ,         �����         �     �� ���       ���� � ������������s          ����	              0   0         �����  L       �     �� ���       ���� � ������������s          ����	              4   4         �����  �       �     �� ���       ���� � ������������s          ����	              8   8         �����  �       �     �� ���       ���� � ������������s          ����	              <   <         ����           �     �� ���       ���� � ������������s          ����	              @   @         ����  <       �	     �� ���       ���� � ������������s          ����	              .  .         �����  �.       �      �� ���        ���� � ������������t          ����	              2  2         �����  v/       �     �� ���        ���� � ������������t          ����	  	 
           6  6         ����  *0       �     �� ���        ���� � ������������t          ����	              :  :         ����J  �0       �     �� ���       ���� � ������������t          ����	              >  >         �����  �1       �     �� ���       ���� � ������������t          ����	              B  B         �����  F2       �     �� ���       ���� � ������������t          ����	              F  F         �����  �2       �     �� ���       ���� � ������������t          ����	              J ! J         ����:  �3       �     �� ���       ���� � ������������t          ����	              N # N         ����v  b4       �     �� ���       ���� � ������������t          ����	              R % R         �����  5       �	     �� ���       ���� � ������������t         ����	  	 
           ?  ?        �����  �J       �      �� ���        ���� � ������������u         ����	              D  D        �����  �K       �     �� ���        ���� � ������������u         ����	              I  I        ����V  XM       �     �� ���        ���� � ������������u         ����	              N  N        �����  �N       �     �� ���       ���� � ������������u         ����	              S  S        ����
  (P       �     �� ���       ���� � ������������u         ����	              X   X "       ����d  �Q       �     �� ���       ���� � ������������u         ����	              ] # ] %       �����  �R       �     �� ���       ���� � ������������u         ����	              b & b (       ����  `T       �     �� ���       ���� � ������������u         ����	              g ) g +       ����r  �U       �     �� ���       ���� � ������������u         ����	              l , l .       �����  0W       �	     �� ���       ���� � ������������u         ����	              Y  Y        ����4  t       �      �� ���        ���� � ������������v         ����	              ^  ^        �����  \v       �     �� ���        ���� � ������������v         ����	              c  c !       ����$  �x       �     �� ���        ���� � ������������v         ����	              h " h $       �����  {       �     �� ���       ���� � ������������v         ����	              m % m '       ����  d}       �     �� ���       ���� � ������������v         ����	              r ( r *       �����  �       �     �� ���       ���� � ������������v         ����	              w + w -       ����  �       �     �� ���       ���� � ������������v         ����	              | . | 0       ����|  l�       �     �� ���       ���� � ������������v         ����	              � 1 � 3       �����  Ć       �     �� ���       ���� � ������������v         ����	    !           � 4 � 6       ����l  �       �	     �� ���       ���� � ������������v         ����	              r   r "       ����L  ȯ       �      �� ���        ���� � ������������w         ����	              w # w %       �����  L�       �     �� ���        ���� � ������������w         ����	              | & | (       ����x  ж       �     �� ���        ���� � ������������w         ����	              � ) � +       ����  T�       �     �� ���       ���� � ������������w         ����	              � , � .       �����  ؽ       �     �� ���       ���� � ������������w         ����	              � / � 1       ����:   \�       �     �� ���       ���� � ������������w         ����	              � 2 � 4       �����   ��       �     �� ���       ���� � ������������w         ����	    !           � 5 � 7       ����f!  d�       �     �� ���       ���� � ������������w         ����	  " #           � 8 � :       �����!  ��    
   �     �� ���       ���� � ������������w         ����	  $ %           � ; � =       �����"  l�    	   �	     �� ���       ���� � ������������w         ����	              � ' � )       �����$  f             �� ���        ���� � ������������x         ����	              � * � ,       �����%  R            �� ���        ���� � ������������x         ����	              � - � /       ����R&  >            �� ���        ���� � ������������x         ����	              � 0 � 2       ����'  *            �� ���       ���� � ������������x         ����	              � 3 � 5       �����'              �� ���       ���� � ������������x         ����	    !           � 6 � 8       ����n(              �� ���       ���� � ������������x         ����	  " #           � 9 � ;       ����")  �            �� ���       ���� � ������������x         ����	  $ %           � < � >       �����)  �$   	         �� ���       ���� � ������������x         ����	  & '           � ? � A       �����*  �)            �� ���       ���� � ������������x         ����	  ( )           � B � D       ����>+  �.       	     �� ���       ���� � ������������x         ����	              � - � /       ����.  pp            �� ���        ���� � �����  �  y         ����	              � 1 � 3       �����.   w           �� ���        ���� � �����  �  y         ����	              � 5 � 7       �����/  �}           �� ���        ���� � �����  �  y         ����	               � 9 � ;       �����0   �           �� ���       ���� � �����  �  y         ����	  ! "           � = � ?       ����V1  ��           �� ���       ���� � �����  �  y         ����	  $ %           � A � C       ����(2  @�   	        �� ���       ���� � �����  �  y         ����	  & '           � E � G       �����2  З           �� ���       ���� � �����  �  y         ����	  ( )           � I � K       �����3  `�           �� ���       ���� � �����  �  y         ����	  * +           � M � O       �����4  �           �� ���       ���� � �����  �  y         ����	  , -           � Q � S       ����p5  ��      	     �� ���       ���� � �����  �  y         ����	              � = � ?       �����8  x�            �� ���        ���� � �����  �  z         ����	               � A � C       �����9  �           �� ���        ���� � �����  �  z         ����	  ! "           � E � G       �����:  X           �� ���        ���� � �����  �  z         ����	  # $           � I � K       �����;  �   	        �� ���       ���� � �����  �  z         ����	  % &           � M � O       ����x<  8            �� ���       ���� � �����  �  z         ����	  ' (           � Q � S       ����h=  �(           �� ���       ���� � �����  �  z         ����	  * +           � U � W       ����X>  1           �� ���       ���� � �����  �  z         ����	  , -           � Y � [       ����H?  �9           �� ���       ���� � �����  �  z         ����	  . /           � ] � _       ����8@  �A           �� ���       ���� � �����  �  z         ����	  0 1           � a � c       ����(A  hJ      	     �� ���       ���� � �����  �  z         ����	  ! "           � L � N       �����D  �            �� ���        ����	 � �����  �  {         ����	  # $           � P � R       �����E  ��   
        �� ���        ����	 � �����  �  {         ����	  % &           � T � V       ����G  (�           �� ���        ����	 � �����  �  {         ����	  ' (           � X � Z       ����H  ��           �� ���       ����	 � �����  �  {         ����	  ) *           � \ � ^       ���� I  @�           �� ���       ����	 � �����  �  {         ����	  + ,           ` b       ����.J  ��           �� ���       ����	 � �����  �  {         ����	  . /           d f       ����<K  X�           �� ���       ����	 � �����  �  {         ����	  0 1           h j       ����JL  ��           �� ���       ����	 � �����  �  {         ����	  2 3           l n       ����XM  p            �� ���       ����	 � �����  �  {         ����	  4 5           p r       ����fN  �   ��  	     �� ���       ����	 � �����  �  {         ����
              � T - !       �����  h�       ;      �� ���        ���� � ������������|         ����
              � X 0 $       ����R  �       ;     �� ���        ���� � ������������|         ����
              � \ 3 '       �����  p�       ;     �� ���        ���� � ������������|         ����
               � ` 6 *       ����~  ��       ;     �� ���       ���� � ������������|         ����
  ! "           � d 9 -       ����  x�       ;     �� ���       ���� � ������������|         ����
  # $           � h < 0       �����  ��       ;     �� ���       ���� � ������������|         ����
  % &           � l ? 3       ����@  ��       ;     �� ���       ���� � ������������|         ����
  ' (           � p B 6       �����  �       ;     �� ���       ���� � ������������|         ����
  * +           � t E 9       ����l   ��    
   ;     �� ���       ���� � ������������|         ����
  , -           � x H <       ����!  �    	   ;	     �� ���       ���� � ������������|         ����
              � c 4 (       ����Z#  v�       <      �� ���        ���� � ������������}         ����
               � h 7 +       ����$  b�       <     �� ���        ���� � ������������}         ����
  ! "           � m : .       �����$  N      <     �� ���        ���� � ������������}         ����
  $ %           � r = 1       ����v%  :      <     �� ���       ���� � ������������}         ����
  & '           � w @ 4       ����*&  &      <     �� ���       ���� � ������������}         ����
  ( )           � | C 7       �����&        <     �� ���       ���� � ������������}         ����
  * +           � � F :       �����'  �      <     �� ���       ���� � ������������}         ����
  , -           � � I =       ����F(  �   	   <     �� ���       ���� � ������������}         ����
  / 0           � � L @       �����(  �      <     �� ���       ���� � ������������}         ����
  1 2           � � O C       �����)  �#      <	     �� ���       ���� � ������������}         ����
  " #           � { : .       ����~,  �c      =      �� ���        ���� � �����  �  ~         ����
  $ %           � � > 2       ����P-  �j      =     �� ���        ���� � �����  �  ~         ����
  & '           � � B 6       ����".  q      =     �� ���        ���� � �����  �  ~         ����
  ) *           � � F :       �����.  �w      =     �� ���       ���� � �����  �  ~         ����
  + ,           � � J >       �����/  0~      =     �� ���       ���� � �����  �  ~         ����
  - .           � N B       �����0  ��   	   =     �� ���       ���� � �����  �  ~         ����
  / 0           � R F       ����j1  P�      =     �� ���       ���� � �����  �  ~         ����
  1 2           � V J       ����<2  ��      =     �� ���       ���� � �����  �  ~         ����
  4 5           � Z N       ����3  p�      =     �� ���       ���� � �����  �  ~         ����
  6 7           � ^ R       �����3   �      =	     �� ���       ���� � �����  �  ~         ����
  ' (           � J >       ����(7  h�      >      �� ���        ���� � �����  �           ����
  ) *           � N B       ����8  ��      >     �� ���        ���� � �����  �           ����
  + ,           � R F       ����9  H      >     �� ���        ���� � �����  �           ����
  . /           � V J       �����9  �	   	   >     �� ���       ���� � �����  �           ����
  0 1            � Z N       �����:  (      >     �� ���       ���� � �����  �           ����
  2 3           '� ^ R       �����;  �      >     �� ���       ���� � �����  �           ����
  4 5           .� b V       �����<  #      >     �� ���       ���� � �����  �           ����
  6 7           5� f Z       �����=  x+      >     �� ���       ���� � �����  �           ����
  9 :           <� j ^       �����>  �3      >     �� ���       ���� � �����  �           ����
  ; <           C� n b       �����?  X<      >	     �� ���       ���� � �����  �           ����
  , -           -� Y M       ����XC  p�      ?      �� ���        ����	 � �����  �  �         ����
  . /           4� ] Q       ����fD  ��   
   ?     �� ���        ����	 � �����  �  �         ����
  0 1           ;� a U       ����tE  ��      ?     �� ���        ����	 � �����  �  �         ����
  3 4           B� e Y       �����F  �      ?     �� ���       ����	 � �����  �  �         ����
  5 6           I� i ]       �����G  ��      ?     �� ���       ����	 � �����  �  �         ����
  7 8           P� m a       �����H  ,�      ?     �� ���       ����	 � �����  �  �         ����
  9 :           W� q e       �����I  ��      ?     �� ���       ����	 � �����  �  �         ����
  ; <           ^� u i       �����J  D�      ?     �� ���       ����	 � �����  �  �         ����
  > ?           e� y m       �����K  ��       ?     �� ���       ����	 � �����  �  �         ����
  @ A           l� } q       �����L  \    ��  ?	     �� ���       ����	 � �����  �  �         ����
              < Y � '       �����  h�       J      �� ���        ���� � �������������         ����
              ? ] � *       ����R  �       J     �� ���        ���� � �������������         ����
              B a � -       �����  p�       J     �� ���        ���� � �������������         ����
              E e � 0       ����~  ��       J     �� ���       ���� � �������������         ����
              H i � 3       ����  x�       J     �� ���       ���� � �������������         ����
              K m � 6       �����  ��       J     �� ���       ���� � �������������         ����
               N q � 9       ����@  ��       J     �� ���       ���� � �������������         ����
  ! "           Q u � <       �����  �       J     �� ���       ���� � �������������         ����
  # $           T y � ?       ����l   ��    
   J     �� ���       ���� � �������������         ����
  % &           W } � B       ����!  �    	   J	     �� ���       ���� � �������������         ����
              C h � .       ����Z#  v�       K      �� ���        ���� � �������������         ����
              G l � 1       ����$  b�       K     �� ���        ���� � �������������         ����
              K p � 4       �����$  N      K     �� ���        ���� � �������������         ����
              O t � 7       ����v%  :      K     �� ���       ���� � �������������         ����
              S x � :       ����*&  &      K     �� ���       ���� � �������������         ����
  ! "           W | � =       �����&        K     �� ���       ���� � �������������         ����
  # $           [ � � @       �����'  �      K     �� ���       ���� � �������������         ����
  % &           _ � � C       ����F(  �   	   K     �� ���       ���� � �������������         ����
  ' (           c � � F       �����(  �      K     �� ���       ���� � �������������         ����
  ) *           g � � I       �����)  �#      K	     �� ���       ���� � �������������         ����
              S w � 4       ����~,  �c      L      �� ���        ���� � �����  �  �         ����
              W | � 8       ����P-  �j      L     �� ���        ���� � �����  �  �         ����
              [ � � <       ����".  q      L     �� ���        ���� � �����  �  �         ����
    !           _ � � @       �����.  �w      L     �� ���       ���� � �����  �  �         ����
  " #           c � � D       �����/  0~      L     �� ���       ���� � �����  �  �         ����
  $ %           g � � H       �����0  ��   	   L     �� ���       ���� � �����  �  �         ����
  ' (           k � L       ����j1  P�      L     �� ���       ���� � �����  �  �         ����
  ) *           o � P       ����<2  ��      L     �� ���       ���� � �����  �  �         ����
  + ,           s � T       ����3  p�      L     �� ���       ���� � �����  �  �         ����
  - .           w � X       �����3   �      L	     �� ���       ���� � �����  �  �         ����
              c � � D       ����(7  h�      M      �� ���        ���� � �����  �  �         ����
    !           g � H       ����8  ��      M     �� ���        ���� � �����  �  �         ����
  " #           k � L       ����9  H      M     �� ���        ���� � �����  �  �         ����
  $ %           o � P       �����9  �	   	   M     �� ���       ���� � �����  �  �         ����
  & '           s � T       �����:  (      M     �� ���       ���� � �����  �  �         ����
  ( )           w �  X       �����;  �      M     �� ���       ���� � �����  �  �         ����
  + ,           { � '\       �����<  #      M     �� ���       ���� � �����  �  �         ����
  - .            � .`       �����=  x+      M     �� ���       ���� � �����  �  �         ����
  / 0           � � 5d       �����>  �3      M     �� ���       ���� � �����  �  �         ����
  1 2           � � <h       �����?  X<      M	     �� ���       ���� � �����  �  �         ����
  " #           r � &S       ����XC  p�      N      �� ���        ����	 � �����  �  �         ����
  $ %           v � -W       ����fD  ��   
   N     �� ���        ����	 � �����  �  �         ����
  & '           z � 4[       ����tE  ��      N     �� ���        ����	 � �����  �  �         ����
  ( )           ~ � ;_       �����F  �      N     �� ���       ����	 � �����  �  �         ����
  * +           � � Bc       �����G  ��      N     �� ���       ����	 � �����  �  �         ����
  , -           � � Ig       �����H  ,�      N     �� ���       ����	 � �����  �  �         ����
  / 0           � � Pk       �����I  ��      N     �� ���       ����	 � �����  �  �         ����
  1 2           � � Wo       �����J  D�      N     �� ���       ����	 � �����  �  �         ����
  3 4           � � ^s       �����K  ��       N     �� ���       ����	 � �����  �  �         ����
  5 6           � � ew       �����L  \    ��  N	     �� ���       ����	 � �����  �  �          ����
              )   )         �����  t1       U      �� ���        ���� � �������������          ����
              -   -         �����  <       U     �� ���        ���� � �������������          ����
              1   1         �����  x       U     �� ���        ���� � �������������          ����
              5   5         �����  �       U     �� ���       ���� � �������������          ����
  	 
           9   9         �����  �       U     �� ���       ���� � �������������          ����
              =   =         ����  ,       U     �� ���       ���� � �������������          ����
              A   A         ����4  h       U     �� ���       ���� � �������������          ����
              E   E         ����R  �       U     �� ���       ���� � �������������          ����
              I   I         ����p  �       U     �� ���       ���� � �������������          ����
              M   M         �����         U	     �� ���       ���� � �������������          ����
              ;  ;         ����  *       V      �� ���        ���� � �������������          ����
              ?  ?         ����B  �*       V     �� ���        ���� � �������������          ����
  	 
           C  C         ����~  z+       V     �� ���        ���� � �������������          ����
              G  G         �����  .,       V     �� ���       ���� � �������������          ����
              K  K         �����  �,       V     �� ���       ���� � �������������          ����
              O  O         ����2  �-       V     �� ���       ���� � �������������          ����
              S  S         ����n  J.       V     �� ���       ���� � �������������          ����
              W ! W         �����  �.       V     �� ���       ���� � �������������          ����
              [ # [         �����  �/       V     �� ���       ���� � �������������          ����
              _ % _         ����"  f0       V	     �� ���       ���� � �������������         ����
  	 
           L  L        ����  HD       W      �� ���        ���� � �������������         ����
              Q  Q        ����l  �E       W     �� ���        ���� � �������������         ����
              V  V        �����  G       W     �� ���        ���� � �������������         ����
              [  [        ����   �H       W     �� ���       ���� � �������������         ����
              `  `        ����z  �I       W     �� ���       ���� � �������������         ����
              e   e "       �����  PK       W     �� ���       ���� � �������������         ����
              j # j %       ����.  �L       W     �� ���       ���� � �������������         ����
              o & o (       �����   N       W     �� ���       ���� � �������������         ����
              t ) t +       �����  �O       W     �� ���       ���� � �������������         ����
              y , y .       ����<  �P       W	     �� ���       ���� � �������������         ����
              f  f        �����  4l       X      �� ���        ���� � �������������         ����
              k  k        ����  �n       X     �� ���        ���� � �������������         ����
              p  p !       �����  �p       X     �� ���        ���� � �������������         ����
              u " u $       ����  <s       X     �� ���       ���� � �������������         ����
              z % z '       �����  �u       X     �� ���       ���� � �������������         ����
               (  *       �����  �w       X     �� ���       ���� � �������������         ����
              � + � -       ����t  Dz       X     �� ���       ���� � �������������         ����
              � . � 0       �����  �|       X     �� ���       ���� � �������������         ����
              � 1 � 3       ����d  �~       X     �� ���       ���� � �������������         ����
    !           � 4 � 6       �����  L�       X	     �� ���       ���� � �������������         ����
                  "       �����  h�       Y      �� ���        ���� � �������������         ����
              � # � %       ����R  �       Y     �� ���        ���� � �������������         ����
              � & � (       �����  p�       Y     �� ���        ���� � �������������         ����
              � ) � +       ����~  ��       Y     �� ���       ���� � �������������         ����
              � , � .       ����  x�       Y     �� ���       ���� � �������������         ����
              � / � 1       �����  ��       Y     �� ���       ���� � �������������         ����
              � 2 � 4       ����@  ��       Y     �� ���       ���� � �������������         ����
    !           � 5 � 7       �����  �       Y     �� ���       ���� � �������������         ����
  " #           � 8 � :       ����l   ��    
   Y     �� ���       ���� � �������������         ����
  $ %           � ; � =       ����!  �    	   Y	     �� ���       ���� � �������������         ����
              � ' � )       ����Z#  v�       Z      �� ���        ���� � �������������         ����
              � * � ,       ����$  b�       Z     �� ���        ���� � �������������         ����
              � - � /       �����$  N      Z     �� ���        ���� � �������������         ����
              � 0 � 2       ����v%  :      Z     �� ���       ���� � �������������         ����
              � 3 � 5       ����*&  &      Z     �� ���       ���� � �������������         ����
    !           � 6 � 8       �����&        Z     �� ���       ���� � �������������         ����
  " #           � 9 � ;       �����'  �      Z     �� ���       ���� � �������������         ����
  $ %           � < � >       ����F(  �   	   Z     �� ���       ���� � �������������         ����
  & '           � ? � A       �����(  �      Z     �� ���       ���� � �������������         ����
  ( )           � B � D       �����)  �#      Z	     �� ���       ���� � �������������         ����
              � - � /       ����~,  �c      [      �� ���        ���� � �����  �  �         ����
              � 1 � 3       ����P-  �j      [     �� ���        ���� � �����  �  �         ����
              � 5 � 7       ����".  q      [     �� ���        ���� � �����  �  �         ����
               � 9 � ;       �����.  �w      [     �� ���       ���� � �����  �  �         ����
  ! "           � = � ?       �����/  0~      [     �� ���       ���� � �����  �  �         ����
  $ %           � A � C       �����0  ��   	   [     �� ���       ���� � �����  �  �         ����
  & '           � E � G       ����j1  P�      [     �� ���       ���� � �����  �  �         ����
  ( )           � I � K       ����<2  ��      [     �� ���       ���� � �����  �  �         ����
  * +           � M � O       ����3  p�      [     �� ���       ���� � �����  �  �         ����
  , -           � Q � S       �����3   �      [	     �� ���       ���� � �����  �  �         ����
              � = � ?       ����(7  h�      \      �� ���        ���� � �����  �  �         ����
               � A � C       ����8  ��      \     �� ���        ���� � �����  �  �         ����
  ! "           � E � G       ����9  H      \     �� ���        ���� � �����  �  �         ����
  # $           � I � K       �����9  �	   	   \     �� ���       ���� � �����  �  �         ����
  % &           � M � O       �����:  (      \     �� ���       ���� � �����  �  �         ����
  ' (           � Q � S       �����;  �      \     �� ���       ���� � �����  �  �         ����
  * +           � U � W       �����<  #      \     �� ���       ���� � �����  �  �         ����
  , -           � Y � [       �����=  x+      \     �� ���       ���� � �����  �  �         ����
  . /           ] _       �����>  �3      \     �� ���       ���� � �����  �  �         ����
  0 1           a c       �����?  X<      \	     �� ���       ���� � �����  �  �         ����
  ! "           � L � N       ����XC  p�      ]      �� ���        ����	 � �����  �  �         ����
  # $           � P � R       ����fD  ��   
   ]     �� ���        ����	 � �����  �  �         ����
  % &           � T � V       ����tE  ��      ]     �� ���        ����	 � �����  �  �         ����
  ' (           X Z       �����F  �      ]     �� ���       ����	 � �����  �  �         ����
  ) *           	\ 	^       �����G  ��      ]     �� ���       ����	 � �����  �  �         ����
  + ,           ` b       �����H  ,�      ]     �� ���       ����	 � �����  �  �         ����
  . /           d f       �����I  ��      ]     �� ���       ����	 � �����  �  �         ����
  0 1           h j       �����J  D�      ]     �� ���       ����	 � �����  �  �         ����
  2 3           !l !n       �����K  ��       ]     �� ���       ����	 � �����  �  �         ����
  4 5           'p 'r       �����L  \    ��  ]	     �� ���       ����	 � �����  �  �         ����              � T - !       ����0   g       �      �� ���        ���� � �������������         ����              � X 0 $       �����  �j       �     �� ���        ���� � �������������         ����              � \ 3 '       ����\  (n       �     �� ���        ���� � �������������         ����    !           � ` 6 *       �����  �q       �     �� ���       ���� � �������������         ����  " #           � d 9 -       �����  0u       �     �� ���       ���� � �������������         ����  $ %           � h < 0       ����  �x       �     �� ���       ���� � �������������         ����  & '           � l ? 3       �����  8|       �     �� ���       ���� � �������������         ����  ( )           � p B 6       ����J  �       �     �� ���       ���� � �������������         ����  + ,           � t E 9       �����  @�    
   �     �� ���       ���� � �������������         ����  - .           � x H <       ����v  Ć    	   �	     �� ���       ���� � �������������         ����              � c 4 (       �����  ��       �      �� ���        ���� � �������������         ����    !           � h 7 +       �����  ��       �     �� ���        ���� � �������������         ����  " #           � m : .       ����6  z�       �     �� ���        ���� � �������������         ����  % &           � r = 1       �����  f�       �     �� ���       ���� � �������������         ����  ' (           � w @ 4       �����  R�       �     �� ���       ���� � �������������         ����  ) *           � | C 7       ����R  >�       �     �� ���       ���� � �������������         ����  + ,           � � F :       ����  *�       �     �� ���       ���� � �������������         ����  - .           � � I =       �����  �    	   �     �� ���       ���� � �������������         ����  0 1            � L @       ����n  �       �     �� ���       ���� � �������������         ����  2 3           � O C       ����"  ��       �	     �� ���       ���� � �������������         ����  # $           � { : .       �����!  �      �      �� ���        ���� � �����  �  �         ����  % &           � � > 2       �����"         �     �� ���        ���� � �����  �  �         ����  ' (           � � B 6       �����#  �      �     �� ���        ���� � �����  �  �         ����  * +           � F :       ����h$  @#      �     �� ���       ���� � �����  �  �         ����  , -           	� J >       ����:%  �)      �     �� ���       ���� � �����  �  �         ����  . /           � N B       ����&  `0   	   �     �� ���       ���� � �����  �  �         ����  0 1           � R F       �����&  �6      �     �� ���       ���� � �����  �  �         ����  2 3           � V J       �����'  �=      �     �� ���       ���� � �����  �  �         ����  5 6           !� Z N       �����(  D      �     �� ���       ���� � �����  �  �         ����  7 8           '� ^ R       ����T)  �J      �	     �� ���       ���� � �����  �  �         ����  ( )           � J >       �����,  |�      �      �� ���        ���� � �����  �  �         ����  * +           � N B       �����-  �      �     �� ���        ���� � �����  �  �         ����  , -           � R F       ����|.  \�      �     �� ���        ���� � �����  �  �         ����  / 0           &� V J       ����l/  ̪   	   �     �� ���       ���� � �����  �  �         ����  1 2           -� Z N       ����\0  <�      �     �� ���       ���� � �����  �  �         ����  3 4           4� ^ R       ����L1  ��      �     �� ���       ���� � �����  �  �         ����  5 6           ;� b V       ����<2  �      �     �� ���       ���� � �����  �  �         ����  7 8           B� f Z       ����,3  ��      �     �� ���       ���� � �����  �  �         ����  : ;           I� j ^       ����4  ��      �     �� ���       ���� � �����  �  �         ����  < =           P� n b       ����5  l�      �	     �� ���       ���� � �����  �  �         ����  - .           :� Y M       �����8  �7      �      �� ���        ����	 � �����  �  �         ����  / 0           A� ] Q       �����9  �B   
   �     �� ���        ����	 � �����  �  �         ����  1 2           H� a U       �����:  M      �     �� ���        ����	 � �����  �  �         ����  4 5           O� e Y       �����;  �W      �     �� ���       ����	 � �����  �  �         ����  6 7           V� i ]       ����=  (b      �     �� ���       ����	 � �����  �  �         ����  8 9           ]� m a       ����>  �l      �     �� ���       ����	 � �����  �  �         ����  : ;           d� q e       ���� ?  @w      �     �� ���       ����	 � �����  �  �         ����  < =           k� u i       ����.@  ́      �     �� ���       ����	 � �����  �  �         ����  ? @           r� y m       ����<A  X�       �     �� ���       ����	 � �����  �  �         ����  A B           y� } q       ����JB  �   ��  �	     �� ���       ����	 � �����  �  �         ����              H f � '       ����0   g       �      �� ���        ���� � �������������         ����              K j � *       �����  �j       �     �� ���        ���� � �������������         ����              N n � -       ����\  (n       �     �� ���        ���� � �������������         ����              Q r � 0       �����  �q       �     �� ���       ���� � �������������         ����              T v � 3       �����  0u       �     �� ���       ���� � �������������         ����              W z � 6       ����  �x       �     �� ���       ���� � �������������         ����    !           Z ~ � 9       �����  8|       �     �� ���       ���� � �������������         ����  " #           ] � � <       ����J  �       �     �� ���       ���� � �������������         ����  $ %           ` � � ?       �����  @�    
   �     �� ���       ���� � �������������         ����  & '           c � � B       ����v  Ć    	   �	     �� ���       ���� � �������������         ����              O u � .       �����  ��       �      �� ���        ���� � �������������         ����              S y � 1       �����  ��       �     �� ���        ���� � �������������         ����              W } � 4       ����6  z�       �     �� ���        ���� � �������������         ����              [ � � 7       �����  f�       �     �� ���       ���� � �������������         ����               _ � � :       �����  R�       �     �� ���       ���� � �������������         ����  " #           c � � =       ����R  >�       �     �� ���       ���� � �������������         ����  $ %           g � � @       ����  *�       �     �� ���       ���� � �������������         ����  & '           k � � C       �����  �    	   �     �� ���       ���� � �������������         ����  ( )           o � � F       ����n  �       �     �� ���       ���� � �������������         ����  * +           s � � I       ����"  ��       �	     �� ���       ���� � �������������         ����              _ � � 4       �����!  �      �      �� ���        ���� � �����  �  �         ����              c � � 8       �����"         �     �� ���        ���� � �����  �  �         ����               g � � <       �����#  �      �     �� ���        ���� � �����  �  �         ����  ! "           k � � @       ����h$  @#      �     �� ���       ���� � �����  �  �         ����  # $           o � D       ����:%  �)      �     �� ���       ���� � �����  �  �         ����  % &           s � H       ����&  `0   	   �     �� ���       ���� � �����  �  �         ����  ( )           w � L       �����&  �6      �     �� ���       ���� � �����  �  �         ����  * +           { � P       �����'  �=      �     �� ���       ���� � �����  �  �         ����  , -            � T       �����(  D      �     �� ���       ���� � �����  �  �         ����  . /           � �  X       ����T)  �J      �	     �� ���       ���� � �����  �  �         ����               o � 
D       �����,  |�      �      �� ���        ���� � �����  �  �         ����  ! "           s � H       �����-  �      �     �� ���        ���� � �����  �  �         ����  # $           w � L       ����|.  \�      �     �� ���        ���� � �����  �  �         ����  % &           { � P       ����l/  ̪   	   �     �� ���       ���� � �����  �  �         ����  ' (            � &T       ����\0  <�      �     �� ���       ���� � �����  �  �         ����  ) *           � � -X       ����L1  ��      �     �� ���       ���� � �����  �  �         ����  , -           � � 4\       ����<2  �      �     �� ���       ���� � �����  �  �         ����  . /           � � ;`       ����,3  ��      �     �� ���       ���� � �����  �  �         ����  0 1           � � Bd       ����4  ��      �     �� ���       ���� � �����  �  �         ����  2 3           � � Ih       ����5  l�      �	     �� ���       ���� � �����  �  �         ����  # $           ~ � 3S       �����8  �7      �      �� ���        ����	 � �����  �  �         ����  % &           � � :W       �����9  �B   
   �     �� ���        ����	 � �����  �  �         ����  ' (           � � A[       �����:  M      �     �� ���        ����	 � �����  �  �         ����  ) *           � � H_       �����;  �W      �     �� ���       ����	 � �����  �  �         ����  + ,           � � Oc       ����=  (b      �     �� ���       ����	 � �����  �  �         ����  - .           � � Vg       ����>  �l      �     �� ���       ����	 � �����  �  �         ����  0 1           � � ]k       ���� ?  @w      �     �� ���       ����	 � �����  �  �         ����  2 3           � � do       ����.@  ́      �     �� ���       ����	 � �����  �  �         ����  4 5           � � ks       ����<A  X�       �     �� ���       ����	 � �����  �  �         ����  6 7           � � rw       ����JB  �   ��  �	     �� ���       ����	 � �����  �  �          ����              6   6         �����  X       �      �� ���        ���� � �������������          ����              :   :         ����  $       �     �� ���        ���� � �������������          ����              >   >         ����0  `       �     �� ���        ���� � �������������          ����   	           B   B         ����N  �       �     �� ���       ���� � �������������          ����  
            F   F         ����l  �       �     �� ���       ���� � �������������          ����              J   J         �����         �     �� ���       ���� � �������������          ����              N   N         �����  P       �     �� ���       ���� � �������������          ����              R   R         �����  �       �     �� ���       ���� � �������������          ����              V   V         �����  �       �     �� ���       ���� � �������������          ����              Z   Z         ����         �	     �� ���       ���� � �������������          ����              H  H         ����z  n
       �      �� ���        ���� � �������������          ����   	           L  L         �����  "       �     �� ���        ���� � �������������          ����  
            P  P         �����  �       �     �� ���        ���� � �������������          ����              T  T         ����.  �       �     �� ���       ���� � �������������          ����              X  X         ����j  >       �     �� ���       ���� � �������������          ����              \  \         �����  �       �     �� ���       ���� � �������������          ����              `  `         �����  �       �     �� ���       ���� � �������������          ����              d ! d         ����  Z       �     �� ���       ���� � �������������          ����              h # h         ����Z         �     �� ���       ���� � �������������          ����              l % l         �����  �       �	     �� ���       ���� � �������������         ����  
            Y  Y        �����         �      �� ���        ���� � �������������         ����              ^  ^        �����  �       �     �� ���        ���� � �������������         ����              c  c        ����:  �       �     �� ���        ���� � �������������         ����              h  h        �����  P       �     �� ���       ���� � �������������         ����              m  m        �����  �       �     �� ���       ���� � �������������         ����              r   r "       ����H   !       �     �� ���       ���� � �������������         ����              w # w %       �����  �"       �     �� ���       ���� � �������������         ����              | & | (       �����  �#       �     �� ���       ���� � �������������         ����              � ) � +       ����V	  X%       �     �� ���       ���� � �������������         ����              � , � .       �����	  �&       �	     �� ���       ���� � �������������         ����              s  s        ����  x7       �      �� ���        ���� � �������������         ����              x  x        �����  �9       �     �� ���        ���� � �������������         ����              }  } !       ����  (<       �     �� ���        ���� � �������������         ����              � " � $       �����  �>       �     �� ���       ���� � �������������         ����              � % � '       �����  �@       �     �� ���       ���� � �������������         ����              � ( � *       ����p  0C       �     �� ���       ���� � �������������         ����              � + � -       �����  �E       �     �� ���       ���� � �������������         ����              � . � 0       ����`  �G       �     �� ���       ���� � �������������         ����               � 1 � 3       �����  8J       �     �� ���       ���� � �������������         ����  ! "           � 4 � 6       ����P  �L       �	     �� ���       ���� � �������������         ����              �   � "       ����0   g       �      �� ���        ���� � �������������         ����              � # � %       �����  �j       �     �� ���        ���� � �������������         ����              � & � (       ����\  (n       �     �� ���        ���� � �������������         ����              � ) � +       �����  �q       �     �� ���       ���� � �������������         ����              � , � .       �����  0u       �     �� ���       ���� � �������������         ����              � / � 1       ����  �x       �     �� ���       ���� � �������������         ����               � 2 � 4       �����  8|       �     �� ���       ���� � �������������         ����  ! "           � 5 � 7       ����J  �       �     �� ���       ���� � �������������         ����  # $           � 8 � :       �����  @�    
   �     �� ���       ���� � �������������         ����  % &           � ; � =       ����v  Ć    	   �	     �� ���       ���� � �������������         ����              � ' � )       �����  ��       �      �� ���        ���� � �������������         ����              � * � ,       �����  ��       �     �� ���        ���� � �������������         ����              � - � /       ����6  z�       �     �� ���        ���� � �������������         ����              � 0 � 2       �����  f�       �     �� ���       ���� � �������������         ����              � 3 � 5       �����  R�       �     �� ���       ���� � �������������         ����  ! "           � 6 � 8       ����R  >�       �     �� ���       ���� � �������������         ����  # $           � 9 � ;       ����  *�       �     �� ���       ���� � �������������         ����  % &           � < � >       �����  �    	   �     �� ���       ���� � �������������         ����  ' (           � ? � A       ����n  �       �     �� ���       ���� � �������������         ����  ) *           � B � D       ����"  ��       �	     �� ���       ���� � �������������         ����              � - � /       �����!  �      �      �� ���        ���� � �����  �  �         ����              � 1 � 3       �����"         �     �� ���        ���� � �����  �  �         ����              � 5 � 7       �����#  �      �     �� ���        ���� � �����  �  �         ����    !           � 9 � ;       ����h$  @#      �     �� ���       ���� � �����  �  �         ����  " #           � = � ?       ����:%  �)      �     �� ���       ���� � �����  �  �         ����  $ %           � A � C       ����&  `0   	   �     �� ���       ���� � �����  �  �         ����  ' (           � E � G       �����&  �6      �     �� ���       ���� � �����  �  �         ����  ) *           � I � K       �����'  �=      �     �� ���       ���� � �����  �  �         ����  + ,           � M � O       �����(  D      �     �� ���       ���� � �����  �  �         ����  - .           � Q � S       ����T)  �J      �	     �� ���       ���� � �����  �  �         ����              � = � ?       �����,  |�      �      �� ���        ���� � �����  �  �         ����    !           � A � C       �����-  �      �     �� ���        ���� � �����  �  �         ����  " #           � E � G       ����|.  \�      �     �� ���        ���� � �����  �  �         ����  $ %           � I � K       ����l/  ̪   	   �     �� ���       ���� � �����  �  �         ����  & '           � M � O       ����\0  <�      �     �� ���       ���� � �����  �  �         ����  ( )           � Q � S       ����L1  ��      �     �� ���       ���� � �����  �  �         ����  + ,           U W       ����<2  �      �     �� ���       ���� � �����  �  �         ����  - .           Y [       ����,3  ��      �     �� ���       ���� � �����  �  �         ����  / 0           ] _       ����4  ��      �     �� ���       ���� � �����  �  �         ����  1 2           a c       ����5  l�      �	     �� ���       ���� � �����  �  �         ����  " #           � L � N       �����8  �7      �      �� ���        ����	 � �����  �  �         ����  $ %           P R       �����9  �B   
   �     �� ���        ����	 � �����  �  �         ����  & '           
T 
V       �����:  M      �     �� ���        ����	 � �����  �  �         ����  ( )           X Z       �����;  �W      �     �� ���       ����	 � �����  �  �         ����  * +           \ ^       ����=  (b      �     �� ���       ����	 � �����  �  �         ����  , -           ` b       ����>  �l      �     �� ���       ����	 � �����  �  �         ����  / 0           "d "f       ���� ?  @w      �     �� ���       ����	 � �����  �  �         ����  1 2           (h (j       ����.@  ́      �     �� ���       ����	 � �����  �  �         ����  3 4           .l .n       ����<A  X�       �     �� ���       ����	 � �����  �  �         ����  5 6           4p 4r       ����JB  �   ��  �	     �� ���       ����	 � �����  �  �         ����              � T - !       �����  (�       �      �� ���        ���� � �������������         ����              � X 0 $       ����r  ��       �     �� ���        ���� � �������������         ����              � \ 3 '       ����   0�       �     �� ���        ���� � �������������         ����  ! "           � ` 6 *       �����   ��       �     �� ���       ���� � �������������         ����  # $           � d 9 -       ����4!  8�       �     �� ���       ���� � �������������         ����  % &           � h < 0       �����!  ��       �     �� ���       ���� � �������������         ����  ' (           � l ? 3       ����`"  @�       �     �� ���       ���� � �������������         ����  ) *           � p B 6       �����"  ��       �     �� ���       ���� � �������������         ����  , -           � t E 9       �����#  H�    
   �     �� ���       ���� � �������������         ����  . /           � x H <       ����"$  ��    	   �	     �� ���       ���� � �������������         ����               � c 4 (       ����z&  V      �      �� ���        ���� � �������������         ����  ! "           � h 7 +       ����.'  B      �     �� ���        ���� � �������������         ����  # $           � m : .       �����'  .      �     �� ���        ���� � �������������         ����  & '           � r = 1       �����(        �     �� ���       ���� � �������������         ����  ( )           � w @ 4       ����J)  !      �     �� ���       ���� � �������������         ����  * +           � | C 7       �����)  �%      �     �� ���       ���� � �������������         ����  , -           � F :       �����*  �*      �     �� ���       ���� � �������������         ����  . /           � I =       ����f+  �/   	   �     �� ���       ���� � �������������         ����  1 2           � L @       ����,  �4      �     �� ���       ���� � �������������         ����  3 4           � O C       �����,  �9      �	     �� ���       ���� � �������������         ����  $ %           � { : .       �����/  �|      �      �� ���        ���� � �����  �  �         ����  & '           � > 2       ����p0  ��      �     �� ���        ���� � �����  �  �         ����  ( )           
� B 6       ����B1  �      �     �� ���        ���� � �����  �  �         ����  + ,           � F :       ����2  ��      �     �� ���       ���� � �����  �  �         ����  - .           � J >       �����2  0�      �     �� ���       ���� � �����  �  �         ����  / 0           � N B       �����3  ��   	   �     �� ���       ���� � �����  �  �         ����  1 2           "� R F       �����4  P�      �     �� ���       ���� � �����  �  �         ����  3 4           (� V J       ����\5  �      �     �� ���       ���� � �����  �  �         ����  6 7           .� Z N       ����.6  p�      �     �� ���       ���� � �����  �  �         ����  8 9           4� ^ R       ���� 7   �      �	     �� ���       ���� � �����  �  �         ����  ) *           � J >       ����H:  �      �      �� ���        ���� � �����  �  �         ����  + ,           %� N B       ����8;  �      �     �� ���        ���� � �����  �  �         ����  - .           ,� R F       ����(<  h      �     �� ���        ���� � �����  �  �         ����  0 1           3� V J       ����=  �%   	   �     �� ���       ���� � �����  �  �         ����  2 3           :� Z N       ����>  H.      �     �� ���       ���� � �����  �  �         ����  4 5           A� ^ R       �����>  �6      �     �� ���       ���� � �����  �  �         ����  6 7           H� b V       �����?  (?      �     �� ���       ���� � �����  �  �         ����  8 9           O� f Z       �����@  �G      �     �� ���       ���� � �����  �  �         ����  ; <           V� j ^       �����A  P      �     �� ���       ���� � �����  �  �         ����  = >           ]� n b       �����B  xX      �	     �� ���       ���� � �����  �  �         ����  . /           G� Y M       ����xF  ��      �      �� ���        ����	 � �����  �  �         ����  0 1           N� ] Q       �����G  <�   
   �     �� ���        ����	 � �����  �  �         ����  2 3           U� a U       �����H  ��      �     �� ���        ����	 � �����  �  �         ����  5 6           \� e Y       �����I  T�      �     �� ���       ����	 � �����  �  �         ����  7 8           c� i ]       �����J  ��      �     �� ���       ����	 � �����  �  �         ����  9 :           j� m a       �����K  l�      �     �� ���       ����	 � �����  �  �         ����  ; <           q� q e       �����L  ��      �     �� ���       ����	 � �����  �  �         ����  = >           x� u i       �����M  �
      �     �� ���       ����	 � �����  �  �         ����  @ A           � y m       �����N         �     �� ���       ����	 � �����  �  �         ����  B C           �� } q       �����O  �   ��  �	     �� ���       ����	 � �����  �  �         ����              U s � '       �����  (�       �      �� ���        ���� � �������������         ����              X w � *       ����r  ��       �     �� ���        ���� � �������������         ����              [ { � -       ����   0�       �     �� ���        ���� � �������������         ����              ^  � 0       �����   ��       �     �� ���       ���� � �������������         ����              a � � 3       ����4!  8�       �     �� ���       ���� � �������������         ����              d � � 6       �����!  ��       �     �� ���       ���� � �������������         ����    !           g � � 9       ����`"  @�       �     �� ���       ���� � �������������         ����  " #           j � � <       �����"  ��       �     �� ���       ���� � �������������         ����  $ %           m � � ?       �����#  H�    
   �     �� ���       ���� � �������������         ����  & '           p � � B       ����"$  ��    	   �	     �� ���       ���� � �������������         ����              \ � � .       ����z&  V      �      �� ���        ���� � �������������         ����              ` � � 1       ����.'  B      �     �� ���        ���� � �������������         ����              d � � 4       �����'  .      �     �� ���        ���� � �������������         ����              h � � 7       �����(        �     �� ���       ���� � �������������         ����               l � � :       ����J)  !      �     �� ���       ���� � �������������         ����  " #           p � � =       �����)  �%      �     �� ���       ���� � �������������         ����  $ %           t � � @       �����*  �*      �     �� ���       ���� � �������������         ����  & '           x �  C       ����f+  �/   	   �     �� ���       ���� � �������������         ����  ( )           | � F       ����,  �4      �     �� ���       ���� � �������������         ����  * +           � � I       �����,  �9      �	     �� ���       ���� � �������������         ����              l � � 4       �����/  �|             �� ���        ���� � �����  �  �         ����              p � � 8       ����p0  ��            �� ���        ���� � �����  �  �         ����               t � <       ����B1  �            �� ���        ���� � �����  �  �         ����  ! "           x � 	@       ����2  ��            �� ���       ���� � �����  �  �         ����  # $           | � D       �����2  0�            �� ���       ���� � �����  �  �         ����  % &           � � H       �����3  ��   	         �� ���       ���� � �����  �  �         ����  ( )           � � L       �����4  P�            �� ���       ���� � �����  �  �         ����  * +           � � !P       ����\5  �            �� ���       ���� � �����  �  �         ����  , -           � � 'T       ����.6  p�            �� ���       ���� � �����  �  �         ����  . /           � � -X       ���� 7   �       	     �� ���       ���� � �����  �  �         ����               | � D       ����H:  �            �� ���        ���� � �����  �  �         ����  ! "           � � H       ����8;  �           �� ���        ���� � �����  �  �         ����  # $           � � %L       ����(<  h           �� ���        ���� � �����  �  �         ����  % &           � � ,P       ����=  �%   	        �� ���       ���� � �����  �  �         ����  ' (           � � 3T       ����>  H.           �� ���       ���� � �����  �  �         ����  ) *           � � :X       �����>  �6           �� ���       ���� � �����  �  �         ����  , -           � � A\       �����?  (?           �� ���       ���� � �����  �  �         ����  . /           � � H`       �����@  �G           �� ���       ���� � �����  �  �         ����  0 1           � � Od       �����A  P           �� ���       ���� � �����  �  �         ����  2 3           � � Vh       �����B  xX      	     �� ���       ���� � �����  �  �         ����  # $           � � @S       ����xF  ��            �� ���        ����	 � �����  �  �         ����  % &           � � GW       �����G  <�   
        �� ���        ����	 � �����  �  �         ����  ' (           � � N[       �����H  ��           �� ���        ����	 � �����  �  �         ����  ) *           � � U_       �����I  T�           �� ���       ����	 � �����  �  �         ����  + ,           � � \c       �����J  ��           �� ���       ����	 � �����  �  �         ����  - .           � � cg       �����K  l�           �� ���       ����	 � �����  �  �         ����  0 1           � � jk       �����L  ��           �� ���       ����	 � �����  �  �         ����  2 3           � � qo       �����M  �
           �� ���       ����	 � �����  �  �         ����  4 5           � � xs       �����N              �� ���       ����	 � �����  �  �         ����  6 7           � � w       �����O  �   ��  	     �� ���       ����	 � �����  �  �          ����              C   C         �����  �        	      �� ���        ���� � �������������          ����              G   G         �����  |       	     �� ���        ���� � �������������          ����              K   K         �����  �       	     �� ���        ���� � �������������          ����   	           O   O         �����  �       	     �� ���       ���� � �������������          ����  
            S   S         ����  0        	     �� ���       ���� � �������������          ����              W   W         ����6  l        	     �� ���       ���� � �������������          ����              [   [         ����T  �        	     �� ���       ���� � �������������          ����              _   _         ����r  �        	     �� ���       ���� � �������������          ����              c   c         �����   !       	     �� ���       ���� � �������������          ����              g   g         �����  \!       		     �� ���       ���� � �������������          ����              U  U         ����&  r3       
      �� ���        ���� � �������������          ����   	           Y  Y         ����b  &4       
     �� ���        ���� � �������������          ����  
            ]  ]         �����  �4       
     �� ���        ���� � �������������          ����              a  a         �����  �5       
     �� ���       ���� � �������������          ����              e  e         ����  B6       
     �� ���       ���� � �������������          ����              i  i         ����R  �6       
     �� ���       ���� � �������������          ����              m  m         �����  �7       
     �� ���       ���� � �������������          ����              q ! q         �����  ^8       
     �� ���       ���� � �������������          ����              u # u         ����  9       
     �� ���       ���� � �������������          ����              y % y         ����B  �9       
	     �� ���       ���� � �������������         ����  
            f  f        ����2  �P             �� ���        ���� � �������������         ����              k  k        �����  0R            �� ���        ���� � �������������         ����              p  p        �����  �S            �� ���        ���� � �������������         ����              u  u        ����@   U            �� ���       ���� � �������������         ����              z  z        �����  hV            �� ���       ���� � �������������         ����                  "       �����  �W            �� ���       ���� � �������������         ����              � # � %       ����N  8Y            �� ���       ���� � �������������         ����              � & � (       �����  �Z            �� ���       ���� � �������������         ����              � ) � +       ����  \            �� ���       ���� � �������������         ����              � , � .       ����\  p]       	     �� ���       ���� � �������������         ����              �  �        �����  �{             �� ���        ���� � �������������         ����              �  �        ����<  ,~            �� ���        ���� � �������������         ����              �  � !       �����  ��            �� ���        ���� � �������������         ����              � " � $       ����,  ܂            �� ���       ���� � �������������         ����              � % � '       �����  4�            �� ���       ���� � �������������         ����              � ( � *       ����  ��            �� ���       ���� � �������������         ����              � + � -       �����  �            �� ���       ���� � �������������         ����              � . � 0       ����  <�            �� ���       ���� � �������������         ����               � 1 � 3       �����  ��            �� ���       ���� � �������������         ����  ! "           � 4 � 6       �����  �       	     �� ���       ���� � �������������         ����              �   � "       �����  (�             �� ���        ���� � �������������         ����              � # � %       ����r  ��            �� ���        ���� � �������������         ����              � & � (       ����   0�            �� ���        ���� � �������������         ����              � ) � +       �����   ��            �� ���       ���� � �������������         ����              � , � .       ����4!  8�            �� ���       ���� � �������������         ����              � / � 1       �����!  ��            �� ���       ���� � �������������         ����               � 2 � 4       ����`"  @�            �� ���       ���� � �������������         ����  ! "           � 5 � 7       �����"  ��            �� ���       ���� � �������������         ����  # $           � 8 � :       �����#  H�    
        �� ���       ���� � �������������         ����  % &           � ; � =       ����"$  ��    	   	     �� ���       ���� � �������������         ����              � ' � )       ����z&  V            �� ���        ���� � �������������         ����              � * � ,       ����.'  B           �� ���        ���� � �������������         ����              � - � /       �����'  .           �� ���        ���� � �������������         ����              � 0 � 2       �����(             �� ���       ���� � �������������         ����              � 3 � 5       ����J)  !           �� ���       ���� � �������������         ����  ! "           � 6 � 8       �����)  �%           �� ���       ���� � �������������         ����  # $           � 9 � ;       �����*  �*           �� ���       ���� � �������������         ����  % &           � < � >       ����f+  �/   	        �� ���       ���� � �������������         ����  ' (           � ? � A       ����,  �4           �� ���       ���� � �������������         ����  ) *           � B � D       �����,  �9      	     �� ���       ���� � �������������         ����              � - � /       �����/  �|            �� ���        ���� � �����  �  �         ����              � 1 � 3       ����p0  ��           �� ���        ���� � �����  �  �         ����              � 5 � 7       ����B1  �           �� ���        ���� � �����  �  �         ����    !           � 9 � ;       ����2  ��           �� ���       ���� � �����  �  �         ����  " #           � = � ?       �����2  0�           �� ���       ���� � �����  �  �         ����  $ %           � A � C       �����3  ��   	        �� ���       ���� � �����  �  �         ����  ' (           � E � G       �����4  P�           �� ���       ���� � �����  �  �         ����  ) *           � I � K       ����\5  �           �� ���       ���� � �����  �  �         ����  + ,           � M � O       ����.6  p�           �� ���       ���� � �����  �  �         ����  - .            Q  S       ���� 7   �      	     �� ���       ���� � �����  �  �         ����              � = � ?       ����H:  �            �� ���        ���� � �����  �  �         ����    !           � A � C       ����8;  �           �� ���        ���� � �����  �  �         ����  " #           � E � G       ����(<  h           �� ���        ���� � �����  �  �         ����  $ %           � I � K       ����=  �%   	        �� ���       ���� � �����  �  �         ����  & '           M O       ����>  H.           �� ���       ���� � �����  �  �         ����  ( )           	Q 	S       �����>  �6           �� ���       ���� � �����  �  �         ����  + ,           U W       �����?  (?           �� ���       ���� � �����  �  �         ����  - .           Y [       �����@  �G           �� ���       ���� � �����  �  �         ����  / 0           ] _       �����A  P           �� ���       ���� � �����  �  �         ����  1 2           !a !c       �����B  xX      	     �� ���       ���� � �����  �  �         ����  " #           L N       ����xF  ��            �� ���        ����	 � �����  �  �         ����  $ %           P R       �����G  <�   
        �� ���        ����	 � �����  �  �         ����  & '           T V       �����H  ��           �� ���        ����	 � �����  �  �         ����  ( )           X Z       �����I  T�           �� ���       ����	 � �����  �  �         ����  * +           #\ #^       �����J  ��           �� ���       ����	 � �����  �  �         ����  , -           )` )b       �����K  l�           �� ���       ����	 � �����  �  �         ����  / 0           /d /f       �����L  ��           �� ���       ����	 � �����  �  �         ����  1 2           5h 5j       �����M  �
           �� ���       ����	 � �����  �  �         ����  3 4           ;l ;n       �����N              �� ���       ����	 � �����  �  �         ����  5 6           Ap Ar       �����O  �   ��  	     �� ���       ����	 � �����  �  �         ����              � T - !       ����l   ��       I      �� ���        ���� � �������������         ����              � X 0 $       ����!  �       I     �� ���        ���� � �������������         ����              � \ 3 '       �����!  ��       I     �� ���        ���� � �������������         ����  ! "           � ` 6 *       ����."  �       I     �� ���       ���� � �������������         ����  # $           � d 9 -       �����"  ��       I     �� ���       ���� � �������������         ����  % &           � h < 0       ����Z#  �       I     �� ���       ���� � �������������         ����  ' (           � l ? 3       �����#  ��       I     �� ���       ���� � �������������         ����  ) *           � p B 6       �����$  $�       I     �� ���       ���� � �������������         ����  , -           � t E 9       ����%  ��    
   I     �� ���       ���� � �������������         ����  . /           � x H <       �����%  ,�    	   I	     �� ���       ���� � �������������         ����               � c 4 (       ����
(  F      J      �� ���        ���� � �������������         ����  ! "           � h 7 +       �����(  2      J     �� ���        ���� � �������������         ����  # $           � m : .       ����r)  "      J     �� ���        ���� � �������������         ����  & '           � r = 1       ����&*  
'      J     �� ���       ���� � �������������         ����  ( )           � w @ 4       �����*  �+      J     �� ���       ���� � �������������         ����  * +           � | C 7       �����+  �0      J     �� ���       ���� � �������������         ����  , -           � F :       ����B,  �5      J     �� ���       ���� � �������������         ����  . /           
� I =       �����,  �:   	   J     �� ���       ���� � �������������         ����  1 2           � L @       �����-  �?      J     �� ���       ���� � �������������         ����  3 4           � O C       ����^.  �D      J	     �� ���       ���� � �������������         ����  $ %           { : .       ����.1  p�      K      �� ���        ���� � �����  �  �         ����  & '           � > 2       ���� 2   �      K     �� ���        ���� � �����  �  �         ����  ( )           � B 6       �����2  ��      K     �� ���        ���� � �����  �  �         ����  + ,           � F :       �����3   �      K     �� ���       ���� � �����  �  �         ����  - .           � J >       ����v4  ��      K     �� ���       ���� � �����  �  �         ����  / 0           � N B       ����H5  @�   	   K     �� ���       ���� � �����  �  �         ����  1 2           %� R F       ����6  а      K     �� ���       ���� � �����  �  �         ����  3 4           +� V J       �����6  `�      K     �� ���       ���� � �����  �  �         ����  6 7           1� Z N       �����7  �      K     �� ���       ���� � �����  �  �         ����  8 9           7� ^ R       �����8  ��      K	     �� ���       ���� � �����  �  �         ����  ) *           !� J >       �����;  �      L      �� ���        ���� � �����  �  �         ����  + ,           (� N B       �����<  #      L     �� ���        ���� � �����  �  �         ����  - .           /� R F       �����=  x+      L     �� ���        ���� � �����  �  �         ����  0 1           6� V J       �����>  �3   	   L     �� ���       ���� � �����  �  �         ����  2 3           =� Z N       �����?  X<      L     �� ���       ���� � �����  �  �         ����  4 5           D� ^ R       �����@  �D      L     �� ���       ���� � �����  �  �         ����  6 7           K� b V       ����xA  8M      L     �� ���       ���� � �����  �  �         ����  8 9           R� f Z       ����hB  �U      L     �� ���       ���� � �����  �  �         ����  ; <           Y� j ^       ����XC  ^      L     �� ���       ���� � �����  �  �         ����  = >           `� n b       ����HD  �f      L	     �� ���       ���� � �����  �  �         ����  . /           J� Y M       ����H  P�      M      �� ���        ����	 � �����  �  �         ����  0 1           Q� ] Q       ����I  ��   
   M     �� ���        ����	 � �����  �  �         ����  2 3           X� a U       ����$J  h�      M     �� ���        ����	 � �����  �  �         ����  5 6           _� e Y       ����2K  ��      M     �� ���       ����	 � �����  �  �         ����  7 8           f� i ]       ����@L  ��      M     �� ���       ����	 � �����  �  �         ����  9 :           m� m a       ����NM        M     �� ���       ����	 � �����  �  �         ����  ; <           t� q e       ����\N  �      M     �� ���       ����	 � �����  �  �         ����  = >           {� u i       ����jO  $      M     �� ���       ����	 � �����  �  �         ����  @ A           �� y m       ����xP  �$       M     �� ���       ����	 � �����  �  �         ����  B C           �� } q       �����Q  </   ��  M	     �� ���       ����	 � �����  �  �         ����              X v � '       ����l   ��       X      �� ���        ���� � �������������         ����              [ z � *       ����!  �       X     �� ���        ���� � �������������         ����              ^ ~ � -       �����!  ��       X     �� ���        ���� � �������������         ����              a � � 0       ����."  �       X     �� ���       ���� � �������������         ����              d � � 3       �����"  ��       X     �� ���       ���� � �������������         ����              g � � 6       ����Z#  �       X     �� ���       ���� � �������������         ����    !           j � � 9       �����#  ��       X     �� ���       ���� � �������������         ����  " #           m � � <       �����$  $�       X     �� ���       ���� � �������������         ����  $ %           p � � ?       ����%  ��    
   X     �� ���       ���� � �������������         ����  & '           s � � B       �����%  ,�    	   X	     �� ���       ���� � �������������         ����              _ � � .       ����
(  F      Y      �� ���        ���� � �������������         ����              c � � 1       �����(  2      Y     �� ���        ���� � �������������         ����              g � � 4       ����r)  "      Y     �� ���        ���� � �������������         ����              k � � 7       ����&*  
'      Y     �� ���       ���� � �������������         ����               o � � :       �����*  �+      Y     �� ���       ���� � �������������         ����  " #           s � � =       �����+  �0      Y     �� ���       ���� � �������������         ����  $ %           w � � @       ����B,  �5      Y     �� ���       ���� � �������������         ����  & '           { � C       �����,  �:   	   Y     �� ���       ���� � �������������         ����  ( )            � 	F       �����-  �?      Y     �� ���       ���� � �������������         ����  * +           � � I       ����^.  �D      Y	     �� ���       ���� � �������������         ����              o � � 4       ����.1  p�      Z      �� ���        ���� � �����  �  �         ����              s �  8       ���� 2   �      Z     �� ���        ���� � �����  �  �         ����               w � <       �����2  ��      Z     �� ���        ���� � �����  �  �         ����  ! "           { � @       �����3   �      Z     �� ���       ���� � �����  �  �         ����  # $            � D       ����v4  ��      Z     �� ���       ���� � �����  �  �         ����  % &           � � H       ����H5  @�   	   Z     �� ���       ���� � �����  �  �         ����  ( )           � � L       ����6  а      Z     �� ���       ���� � �����  �  �         ����  * +           � � $P       �����6  `�      Z     �� ���       ���� � �����  �  �         ����  , -           � � *T       �����7  �      Z     �� ���       ���� � �����  �  �         ����  . /           � � 0X       �����8  ��      Z	     �� ���       ���� � �����  �  �         ����                � D       �����;  �      [      �� ���        ���� � �����  �  �         ����  ! "           � � !H       �����<  #      [     �� ���        ���� � �����  �  �         ����  # $           � � (L       �����=  x+      [     �� ���        ���� � �����  �  �         ����  % &           � � /P       �����>  �3   	   [     �� ���       ���� � �����  �  �         ����  ' (           � � 6T       �����?  X<      [     �� ���       ���� � �����  �  �         ����  ) *           � � =X       �����@  �D      [     �� ���       ���� � �����  �  �         ����  , -           � � D\       ����xA  8M      [     �� ���       ���� � �����  �  �         ����  . /           � � K`       ����hB  �U      [     �� ���       ���� � �����  �  �         ����  0 1           � � Rd       ����XC  ^      [     �� ���       ���� � �����  �  �         ����  2 3           � � Yh       ����HD  �f      [	     �� ���       ���� � �����  �  �         ����  # $           � � CS       ����H  P�      \      �� ���        ����	 � �����  �  �         ����  % &           � � JW       ����I  ��   
   \     �� ���        ����	 � �����  �  �         ����  ' (           � � Q[       ����$J  h�      \     �� ���        ����	 � �����  �  �         ����  ) *           � � X_       ����2K  ��      \     �� ���       ����	 � �����  �  �         ����  + ,           � � _c       ����@L  ��      \     �� ���       ����	 � �����  �  �         ����  - .           � � fg       ����NM        \     �� ���       ����	 � �����  �  �         ����  0 1           � � mk       ����\N  �      \     �� ���       ����	 � �����  �  �         ����  2 3           � � to       ����jO  $      \     �� ���       ����	 � �����  �  �         ����  4 5           � � {s       ����xP  �$       \     �� ���       ����	 � �����  �  �         ����  6 7           � � �w       �����Q  </   ��  \	     �� ���       ����	 � �����  �  �          ����              F   F         ����0  �        c      �� ���        ���� � �������������          ����              J   J         ����N  �"       c     �� ���        ���� � �������������          ����              N   N         ����l  �"       c     �� ���        ���� � �������������          ����   	           R   R         �����  #       c     �� ���       ���� � �������������          ����  
            V   V         �����  P#       c     �� ���       ���� � �������������          ����              Z   Z         �����  �#       c     �� ���       ���� � �������������          ����              ^   ^         �����  �#       c     �� ���       ���� � �������������          ����              b   b         ����  $       c     �� ���       ���� � �������������          ����              f   f         ����   @$       c     �� ���       ���� � �������������          ����              j   j         ����>  |$       c	     �� ���       ���� � �������������          ����              X  X         �����  "8       d      �� ���        ���� � �������������          ����   	           \  \         �����  �8       d     �� ���        ���� � �������������          ����  
            `  `         ����.  �9       d     �� ���        ���� � �������������          ����              d  d         ����j  >:       d     �� ���       ���� � �������������          ����              h  h         �����  �:       d     �� ���       ���� � �������������          ����              l  l         �����  �;       d     �� ���       ���� � �������������          ����              p  p         ����  Z<       d     �� ���       ���� � �������������          ����              t ! t         ����Z  =       d     �� ���       ���� � �������������          ����              x # x         �����  �=       d     �� ���       ���� � �������������          ����              | % |         �����  v>       d	     �� ���       ���� � �������������         ����  
            i  i        �����  W       e      �� ���        ���� � �������������         ����              n  n        ����  pX       e     �� ���        ���� � �������������         ����              s  s        ����v  �Y       e     �� ���        ���� � �������������         ����              x  x        �����  @[       e     �� ���       ���� � �������������         ����              }  }        ����*  �\       e     �� ���       ���� � �������������         ����              �   � "       �����  ^       e     �� ���       ���� � �������������         ����              � # � %       �����  x_       e     �� ���       ���� � �������������         ����              � & � (       ����8  �`       e     �� ���       ���� � �������������         ����              � ) � +       �����  Hb       e     �� ���       ���� � �������������         ����              � , � .       �����  �c       e	     �� ���       ���� � �������������         ����              �  �        ����T  ��       f      �� ���        ���� � �������������         ����              �  �        �����  ��       f     �� ���        ���� � �������������         ����              �  � !       ����D  T�       f     �� ���        ���� � �������������         ����              � " � $       �����  ��       f     �� ���       ���� � �������������         ����              � % � '       ����4  �       f     �� ���       ���� � �������������         ����              � ( � *       �����  \�       f     �� ���       ���� � �������������         ����              � + � -       ����$  ��       f     �� ���       ���� � �������������         ����              � . � 0       �����  �       f     �� ���       ���� � �������������         ����               � 1 � 3       ����  d�       f     �� ���       ���� � �������������         ����  ! "           � 4 � 6       �����  ��       f	     �� ���       ���� � �������������         ����              �   � "       ����l   ��       g      �� ���        ���� � �������������         ����              � # � %       ����!  �       g     �� ���        ���� � �������������         ����              � & � (       �����!  ��       g     �� ���        ���� � �������������         ����              � ) � +       ����."  �       g     �� ���       ���� � �������������         ����              � , � .       �����"  ��       g     �� ���       ���� � �������������         ����              � / � 1       ����Z#  �       g     �� ���       ���� � �������������         ����               � 2 � 4       �����#  ��       g     �� ���       ���� � �������������         ����  ! "           � 5 � 7       �����$  $�       g     �� ���       ���� � �������������         ����  # $           � 8 � :       ����%  ��    
   g     �� ���       ���� � �������������         ����  % &           � ; � =       �����%  ,�    	   g	     �� ���       ���� � �������������         ����              � ' � )       ����
(  F      h      �� ���        ���� � �������������         ����              � * � ,       �����(  2      h     �� ���        ���� � �������������         ����              � - � /       ����r)  "      h     �� ���        ���� � �������������         ����              � 0 � 2       ����&*  
'      h     �� ���       ���� � �������������         ����              � 3 � 5       �����*  �+      h     �� ���       ���� � �������������         ����  ! "           � 6 � 8       �����+  �0      h     �� ���       ���� � �������������         ����  # $           � 9 � ;       ����B,  �5      h     �� ���       ���� � �������������         ����  % &           � < � >       �����,  �:   	   h     �� ���       ���� � �������������         ����  ' (           � ? � A       �����-  �?      h     �� ���       ���� � �������������         ����  ) *           � B � D       ����^.  �D      h	     �� ���       ���� � �������������         ����              � - � /       ����.1  p�      i      �� ���        ���� � �����  �  �         ����              � 1 � 3       ���� 2   �      i     �� ���        ���� � �����  �  �         ����              � 5 � 7       �����2  ��      i     �� ���        ���� � �����  �  �         ����    !           � 9 � ;       �����3   �      i     �� ���       ���� � �����  �  �         ����  " #           � = � ?       ����v4  ��      i     �� ���       ���� � �����  �  �         ����  $ %           � A � C       ����H5  @�   	   i     �� ���       ���� � �����  �  �         ����  ' (           � E � G       ����6  а      i     �� ���       ���� � �����  �  �         ����  ) *           � I � K       �����6  `�      i     �� ���       ���� � �����  �  �         ����  + ,           � M � O       �����7  �      i     �� ���       ���� � �����  �  �         ����  - .           Q S       �����8  ��      i	     �� ���       ���� � �����  �  �         ����              � = � ?       �����;  �      j      �� ���        ���� � �����  �  �         ����    !           � A � C       �����<  #      j     �� ���        ���� � �����  �  �         ����  " #           � E � G       �����=  x+      j     �� ���        ���� � �����  �  �         ����  $ %            I  K       �����>  �3   	   j     �� ���       ���� � �����  �  �         ����  & '           M O       �����?  X<      j     �� ���       ���� � �����  �  �         ����  ( )           Q S       �����@  �D      j     �� ���       ���� � �����  �  �         ����  + ,           U W       ����xA  8M      j     �� ���       ���� � �����  �  �         ����  - .           Y [       ����hB  �U      j     �� ���       ���� � �����  �  �         ����  / 0           ] _       ����XC  ^      j     �� ���       ���� � �����  �  �         ����  1 2           $a $c       ����HD  �f      j	     �� ���       ���� � �����  �  �         ����  " #           L N       ����H  P�      k      �� ���        ����	 � �����  �  �         ����  $ %           P R       ����I  ��   
   k     �� ���        ����	 � �����  �  �         ����  & '           T V       ����$J  h�      k     �� ���        ����	 � �����  �  �         ����  ( )            X  Z       ����2K  ��      k     �� ���       ����	 � �����  �  �         ����  * +           &\ &^       ����@L  ��      k     �� ���       ����	 � �����  �  �         ����  , -           ,` ,b       ����NM        k     �� ���       ����	 � �����  �  �         ����  / 0           2d 2f       ����\N  �      k     �� ���       ����	 � �����  �  �         ����  1 2           8h 8j       ����jO  $      k     �� ���       ����	 � �����  �  �         ����  3 4           >l >n       ����xP  �$       k     �� ���       ����	 � �����  �  �         ����  5 6           Dp Dr       �����Q  </   ��  k	     �� ���       ����	 � �����  �  �           g                � � s b       �����?  }       �      ��$ ���        ����   ����������������         g                � � � r       �����I  �O       �      ��$ ���        ����   ����������������         g                � � � �       ����T  A       �      ��$ ���        ����   ����������������         g                
� �       ����A_  QS       �      ��$ ���        ����   ����������������         g                @#� �       ����$k  ��       �      ��$ ��         ����   ����������������         g                m<� �       �����w  ��       �      ��$ ��        ����   ����������������         g                �U� �       �����  <d
       �      ��$ ��        ����   ����������������         g                �s� 	      ������  �       �      ��$ ��        ����   ����������������         g                �'      ������  ��       �      ��$ ��        ����   ����������������         g                :�E      �����  p�       �      ��$ ��        ����   ����������������         g                v�6c      ����%�  x       �      ��$ ��        ����   ����������������        # g                � � � b       �����?  }       �      ��% ��        ����   ����������������        $ g                � � m       �����I  �O       �      ��% ��        ����   ����������������        % g                � � -�       ����T  A       �      ��% ��	        ����   ����������������        & g                P�       ����A_  QS       �      ��% ��
        ����   ����������������        ' g                ?x�       ����$k  ��       �      ��% ��        ����   ����������������        ( g                ,b��       �����w  ��       �      ��% ��        ����   ����������������        ) g                B���       �����  <d
       �      ��% ��        ����   ����������������        * g                W��       ������  �       �      ��% ��        ����   ����������������        + g                k�J�       ������  ��       �      ��% ��        ����   ����������������        , g                ��      �����  p�       �      ��% ��        ����   ����������������        - g                � �$      ����%�  x       �      ��% ��        ����   ����������������          g                            �����   �        �      ��& ��        ����   ����������������        . g                           ����B  �        �      ��& ��        ����   ����������������        / g                          ����[  l        �      ��& ��        ����   ����������������        0 g                &          ����'  �#        �      ��& ��        ����   ����������������        1 g                .  %        �����
  �?        �      ��& ��        ����   ����������������        2 g                A " 6 "       �����  �g        �      ��& ��        ����   ����������������        3 g                L ) @ )       �����  �        �      ��& ��        ����   ����������������        4 g                e 1 W 1       ����U  ��        �      ��& ��        ����   ����������������        5 g                s : d :       �����  @<       �      ��& ��        ����	   ����������������        6 g                � A � A       �����&  ʨ       �      ��& ��        ����
   ����������������        7 g                � L � L       ����O.  �+       �      ��& ��        ����   ����������������        8 g                � U � U       �����6  �       �      ��& ��        ����   ����������������        9 g                � b � b       �����?  }       �      ��& ��        ����   ����������������        : g                � m � m       �����I  �O       �      ��& ��        ����   ����������������        ; g                � �       ����T  A       �      ��& ��         ����   ����������������        < g                ;� )�       ����A_  QS              ��& ��!        ����   ����������������        = g                U� C�       ����$k  ��             ��& ��"        ����   ����������������        > g                q� p�       �����w  ��             ��& ��#        ����   ����������������        ? g                �� ��       �����  <d
             ��& ��$        ����   ����������������        @ g                �"�      ������  �             ��& ��%        ����   ����������������        A g                �J�D      ������  ��             ��& ��&        ����   ����������������        B g                �t.l      �����  p�             ��& ��'        ����   ����������������        C g                ��`�      ����%�  x             ��& ��(        ����   ����������������        ��j ��          2                �����   �              ��@ ��)        ������  ����������������        ��j ��          2                ����B  �              ��A ��*        ������  ����������������        ��j ��          2                ����[  l        	      ��B ��+        ������  ����������������        ����k ��"1                          �����   �        �      ��; ��,        ������  ����������������        ����k ��#1                          �����  �        �      ��; ��-        ������  ����������������        ����k ��$1                          ����  @        �      ��; ��.        ������  ����������������        ����k ��%1                          �����  L"        �      ��; ��/        ������  ����������������        ����k ��&1                          ����r  ��        �      ��< ��0        ������  ����������������        ����k ��'1                          ����
  Z�        �      ��< ��1        ������  ����������������        ����k ��(1                          ����U  R9       �      ��< ��2        ������  ����������������        ����k ��)1                          ����S&  ��       �      ��< ��3        ������  ����������������         ��l ��U        2                  �����   �        �      ��= ��4        ������  ����������������         ��i ��                            �����  C        S     ��6 ��5        ������  ����������������        ����h ��                           �      ]               ��? ��6        ������  ����������������        ����h ��         2                  �                     ��? ��7        ������  ����������������        ����h ��         d                  �      �              ��? ��8        ������  ����������������        ����h ��         �                  �      �              ��? ��9        ������  ����������������        ����h ��         �                  �      n              ��? ��:        ������  ����������������        ����h ��         �                  �      6              ��? ��;        ������  ����������������         ��d ��                         �   �   �        �     ��. ��<        ������  ����������������         ��d ��                         �   �  S        �     ��. ��=        ������  ����������������         ��d ��  (        
               �   �  �        �     ��. ��>        ������  ����������������         ��d ��  2                       �   !  �        �     ��. ��?        ������  ����������������         ��e ��                         �   �   �        �     ��/ ��@        ������  ����������������         ��e ��                         �   �  S        �     ��/ ��A        ������  ����������������         ��e ��  (        
               �   �  �        �     ��/ ��B        ������  ����������������         ��e ��  2                       �   !  �        �     ��/ ��C        ������  ����������������        ��m ��                          P  �   �              ��C ��D        ������  ����������������        ��m ��                          8J  �                ��D ��E        ������  ����������������        ��m ��                          Hq  �  �              ��E ��F        ������  ����������������        ��m ��                         P�    8              ��F ��G        ������  ����������������        ��m ��                         �� �  B'              ��G ��H        ������  ����������������        ��m ��                         @ Y  D              ��H ��I        ������  ����������������        ��m ��                    3     �� �  �l              ��I ��J        ������  ����������������        ��m ��                    L     P� p  ��              ��J ��K        ������  ����������������        ��m ��                    y     ��%   H�              ��K ��L        ������  ����������������          ���3�32    d                �  X                   M    �������c   �������������            ���5�52    i             
     $                  M    �������c   �������������            ���7�72    n                0  `                  M    �������c   �������������            ���9�92    s                N  �                  M   �������c   �������������            ���;�;2    x                l  �                  M   �������c   �������������            ���=�=2    }                �                    M   �������c   �������������            ���?�?2    �                �  P                  M   �������c   �������������            ���A�A2    �                �  �                  M   �������c   �������������            ���C�C2    �                �  �                  M   �������c   �������������            ���E�E2    �                           	         M   �������c   �������������            ��U�R�2        d            �          l       h   N    �������c   �������������            ��W�T�2        i         	   �  �        l      h   N    �������c   �������������            ��Y�V�2        n         
   �  �        l      h   N    �������c   �������������            ��[�X�2        s         
     $        l      h   N   �������c   �������������            ��]�Z�2        x            0  `        l      h   N   �������c   �������������            ��_�\�2        }            N  �        l      h   N   �������c   �������������            ��a�^�2        �            l  �        l      h   N   �������c   �������������            ��c�`�2        �            �          l      h   N   �������c   �������������            ��e�b�2        �            �  P        l      h   N   �������c   �������������            ��g�d�2        �            �  �        l 	     h   N   �������c   �������������             �f�f
2      K K            l  �        �       �   O    Ƭ�����c   �������������             �h�h
2      M O            �          �      �   O    Ƭ�����c   �������������             �j�j
2      O S            �  P        �      �   O    Ƭ�����c   �������������             �l�l
2      Q W            �  �        �      �   O   Ƭ�����c   �������������             �n�n
2      S [            �  �        �      �   O   Ƭ�����c   �������������             �p�p
2      U _                      �      �   O   Ƭ�����c   �������������             �r�r
2      W c               @        �      �   O   Ƭ�����c   �������������             �t�t
2      Y g            >  |        �      �   O   Ƭ�����c   �������������             �v�v
2      [ k            \  �        �      �   O   Ƭ�����c   �������������              x x
2      ] o            z  �        � 	     �   O   Ƭ�����c   �������������         ����� ��                            ����'   N        d      ��P ��P        ������  ����������������       ����� ��                            ����'   N        e      ��P ��Q        ������  ����������������       ����� ��                            ����'   N        f      ��P ��R        ������  ����������������       ����� ��                            ����'   N        g      ��P ��S        ������  ����������������       ����� ��                            ����'   N        h      ��P ��T        ������  ����������������       ����� ��                            ����'   N        i      ��P ��U        ������  ����������������       ����� ��                            ����'   N        j      ��P ��V        ������  ����������������       ����� ��                            ����'   N        k      ��P ��W        ������  ����������������       ����� ��                            ����'   N        l      ��P ��X        ������  ����������������       ����� ��                            ����'   N        m      ��P ��Y        ������  ����������������       ����� ��                            ����'   N        n      ��P ��Z        ������  ����������������       ����� ��                            ����'   N        o      ��P ��[        ������  ����������������       ����� ��                            ����'   N        p      ��P ��\        ������  ����������������       ����� ��                            ����'   N        q      ��P ��]        ������  ����������������       ����� ��                            ����'   N        r      ��P ��^        ������  ����������������       ����� ��                            ����'   N        s      ��P ��_        ������  ����������������       ����� ��                            ����'   N        t      ��P ��`        ������  ����������������       ����� ��                            ����'   N        u      ��P ��a        ������  ����������������       ����� ��                            ����'   N        v      ��P ��b        ������  ����������������       ����� ��                            ����'   N        w      ��P ��c        ������  ����������������       ����� ��                            ����'   N        x      ��P ��d        ������  ����������������       ����� ��                            ����'   N        y      ��P ��e        ������  ����������������       ����� ��                            ����'   N        z      ��P ��f        ������  ����������������       ����� ��                            ����'   N        {      ��P ��g        ������  ����������������       ����� ��                            �����  �        >      ��S ��h        ������  ����������������       ����� ��                            ����'   N        |      ��Q ��i        ������  ����������������       ����� ��                            ����'   N        }      ��Q ��j        ������  ����������������       ����� ��                            ����'   N        ~      ��Q ��k        ������  ����������������       ����� ��                            ����'   N              ��Q ��l        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��m        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��n        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��o        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��p        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��q        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��r        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��s        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��t        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��u        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��v        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��w        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��x        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��y        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��z        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��{        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��|        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��}        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��~        ������  ����������������       ����� ��                            ����'   N        �      ��Q ��        ������  ����������������       ����� ��                            ����'   N        �      ��Q ���        ������  ����������������       ����  < =          � d           2   `	  �        �      �   �        ����c   �������������         ����  > ?          � g           0   ~	  �        �     �   �        ����c   �������������         ����  @ A          � j           1   �	  8        �     �   �        ����c   �������������         ����  B C          � m           1   �	  t        �     �   �       ����c   �������������         ����  D E          � p           2   �	  �        �     �   �       ����c   �������������         ����  F G          � s           3   �	  �        �     �   �       ����c   �������������         ����  H I          � v           3   
  (        �     �   �       ����c   �������������         ����  J K          � y           4   2
  d        �     �   �       ����c   �������������         ����  L M          � |           4   P
  �        �     �   �       ����c   �������������         ����  N O          �            5   n
  �        �	     �   �       ����c   �������������         ����  2 3            d �         2   `	  �        �      �   �        ����c   �������������         ����  4 5            g �         0   ~	  �        �     �   �        ����c   �������������         ����  6 7            j �         1   �	  8        �     �   �        ����c   �������������         ����  8 9            m �         1   �	  t        �     �   �       ����c   �������������         ����  : ;            p �         2   �	  �        �     �   �       ����c   �������������         ����  < =            s �         3   �	  �        �     �   �       ����c   �������������         ����  > ?            v �         3   
  (        �     �   �       ����c   �������������         ����  @ A            y �         4   2
  d        �     �   �       ����c   �������������         ����  B C            | �         4   P
  �        �     �   �       ����c   �������������         ����  D E             �         5   n
  �        �	     �   �       ����c   �������������         ����  1 2          �   �         2   `	  �        �      �   �        ����c   �������������         ����  3 4          �   �         0   ~	  �        �     �   �        ����c   �������������         ����  5 6          �   �         1   �	  8        �     �   �        ����c   �������������         ����  7 8          �   �         1   �	  t        �     �   �       ����c   �������������         ����  9 :          �   �         2   �	  �        �     �   �       ����c   �������������         ����  ; <          �   �         3   �	  �        �     �   �       ����c   �������������         ����  = >          �   �         3   
  (        �     �   �       ����c   �������������         ����  ? @          �   �         4   2
  d        �     �   �       ����c   �������������         ����  A B          �   �         4   P
  �        �     �   �       ����c   �������������         ����  C D          �   �         5   n
  �        �	     �   �       ����c   �������������         ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������        ����               # 1        	      �       R        ���        ���� � �������������          ����               & 6           >  |       R       ���        ���� � �������������          ����               ) ;            \  �       R       ���        ���� � �������������          ����    	           , @ "          z  �       R       ���       ���� � �������������          ����   
            / E $          �  0       R       ���       ���� � �������������          ����                2 J &          �  l       R       ���       ���� � �������������          ����              " 5 O (          �  �       R       ���       ���� � �������������          ����              $ 8 T *          �  �       R       ���       ���� � �������������          ����              & ; Y ,                    R       ���       ���� � �������������          ����              ( > ^ .          .  \       R	       ���       ���� � �������������          ����               + L        #   �  �       S        ���        ���� � �������������          ����               . Q        %   �  �       S       ���        ���� � �������������          ����   	 
           1 V        '     Z       S       ���        ���� � �������������          ����               4 [ !       )   Z         S       ���       ���� � �������������          ����              ! 7 ` #       *   �  �       S       ���       ���� � �������������          ����              $ : e %       ,   �  v       S       ���       ���� � �������������          ����              ' = j '       .     *       S       ���       ���� � �������������          ����              * @ o )       0   J  �       S       ���       ���� � �������������          ����              - C t +       2   �  �       S       ���       ���� � �������������          ����              0 F y -       3   �  F       S	       ���       ���� � �������������          ����    	           2 f        N   �  �       T        ���        ���� � �������������         ����   
             6 k        R     0        T       ���        ���� � �������������         ����              # : p        V   f  �!       T       ���        ���� � �������������         ����              & > u "       Y   �   #       T       ���       ���� � �������������         ����              ) B z %       ]   	  h$       T       ���       ���� � �������������         ����              , F  (       `   t	  �%       T       ���       ���� � �������������         ����              / J � +       d   �	  8'       T       ���       ���� � �������������         ����              2 N � .       h   (
  �(       T       ���       ���� � �������������         ����              5 R � 1       k   �
  *       T       ���       ���� � �������������         ����              8 V � 4       o   �
  p+       T	       ���       ���� � �������������          ����              % C  !       �   D  T=       U        ���        ���� � �������������         ����              ( G � $       �   �  �?       U       ���        ���� � �������������         ����              + K � '       �   4  B       U       ���        ���� � �������������         ����              . O � *       �   �  \D       U       ���       ���� � �������������         ����              1 S � -       �   $  �F       U       ���       ���� � �������������         ����              4 W � 0       �   �  I       U       ���       ���� � �������������         ����              7 [ � 3       �     dK       U       ���       ���� � �������������         ����              : _ � 6       �   �  �M       U       ���       ���� � �������������         ����              = c � 9       �     P       U       ���       ���� � �������������         ����              @ g � <       �   |  lR       U	       ���       ���� � �������������          ����              , S � (         \  (n       V        ���        ���� � �������������         ����              / W � +       #  �  �q       V       ���        ���� � �������������         ����              2 [ � .       ,  �  0u       V       ���        ���� � �������������         ����              5 _ � 1       5    �x       V       ���       ���� � �������������         ����              8 c � 4       >  �  8|       V       ���       ���� � �������������         ����              ; g � 7       G  J  �       V       ���       ���� � �������������         ����              > k � :       P  �  @�       V       ���       ���� � �������������         ����              A o � =       Y  v  Ć       V       ���       ���� � �������������         ����              D s � @       b    H�    
   V       ���       ���� � �������������         ����     !          G w � C       k  �  ̍    	   V	       ���       ���� � �������������          ����               (           ,  h       �        ���        ���� � �������������          ����               -           J  �       �       ���        ���� � �������������          ����                2           h  �       �       ���        ���� � �������������          ����              # 7           �         �       ���       ���� � �������������          ����  	 
           & <           �  H       �       ���       ���� � �������������          ����              ) A        	   �  �       �       ���       ���� � �������������          ����              , F        	   �  �       �       ���       ���� � �������������          ����              / K !       
   �  �       �       ���       ���� � �������������          ����              2 P #       
     8       �       ���       ���� � �������������          ����              5 U %          :  t       �	       ���       ���� � �������������          ����              " C           �         �        ���        ���� � �������������          ����              % H           �  �       �       ���        ���� � �������������          ����   	           ( M           *  ~	       �       ���        ���� � �������������          ����  
            + R           f  2
       �       ���       ���� � �������������          ����              . W           �  �
       �       ���       ���� � �������������          ����              1 \           �  �       �       ���       ���� � �������������          ����              4 a             N       �       ���       ���� � �������������          ����             ! 7 f         !   V         �       ���       ���� � �������������          ����             $ : k "       #   �  �       �       ���       ���� � �������������          ����             ' = p $       $   �  j       �	       ���       ���� � �������������          ����              ) ]        :   �  �       �        ���        ���� � �������������         ����  	 
           - b        >     `       �       ���        ���� � �������������         ����              1 g        B   r  �       �       ���        ���� � �������������         ����              5 l        E   �  0       �       ���       ���� � �������������         ����               9 q        I   &  �       �       ���       ���� � �������������         ����             # = v        L   �          �       ���       ���� � �������������         ����             & A { "       P   �  h       �       ���       ���� � �������������         ����             ) E � %       T   4  �        �       ���       ���� � �������������         ����             , I � (       W   �  8"       �       ���       ���� � �������������         ����             / M � +       [   �  �#       �	       ���       ���� � �������������          ����  
            : v        �   P
  �3       �        ���        ���� � �������������         ����              > |        �   �
  �5       �       ���        ���� � �������������         ����             " B �        �   @  @8       �       ���        ���� � �������������         ����             % F � !       �   �  �:       �       ���       ���� � �������������         ����             ( J � $       �   0  �<       �       ���       ���� � �������������         ����             + N � '       �   �  H?       �       ���       ���� � �������������         ����             . R � *       �      �A       �       ���       ���� � �������������         ����             1 V � -       �   �  �C       �       ���       ���� � �������������         ����             4 Z � 0       �     PF       �       ���       ���� � �������������         ����             7 ^ � 3       �   �  �H       �	       ���       ���� � �������������          ����             # J �        �   h  pb       �        ���        ���� � �������������         ����             & N � "         �  �e       �       ���        ���� � �������������         ����             ) R � %         �  xi       �       ���        ���� � �������������         ����             , V � (         *  �l       �       ���       ���� � �������������         ����             / Z � +          �  �p       �       ���       ���� � �������������         ����             2 ^ � .       )  V  t       �       ���       ���� � �������������         ����             5 b � 1       2  �  �w       �       ���       ���� � �������������         ����             8 f � 4       ;  �  {       �       ���       ���� � �������������         ����             ; j � 7       D    �~    
   �       ���       ���� � �������������         ����              > n � :       M  �  �    	   �	       ���       ���� � �������������          ����              % +           �   �        #        ���        ���� � �������������          ����             ! ( 0           �   �       #       ���        ���� � �������������          ����             # + 5                     #       ���        ���� � �������������          ����             % . : "          "  D       #       ���       ���� � �������������          ����  	 
          ' 1 ? $          @  �       #       ���       ���� � �������������          ����             ) 4 D &          ^  �       #       ���       ���� � �������������          ����             + 7 I (          |  �       #       ���       ���� � �������������          ����             - : N *          �  4       #       ���       ���� � �������������          ����             / = S ,          �  p       #       ���       ���� � �������������          ����             1 @ X .       	   �  �       #	       ���       ���� � �������������          ����              - F           N  �       $        ���        ���� � �������������          ����             ! 0 K           �  �       $       ���        ���� � �������������          ����   	          $ 3 P           �  R       $       ���        ���� � �������������          ����  
           ' 6 U !            	       $       ���       ���� � �������������          ����             * 9 Z #          >  �	       $       ���       ���� � �������������          ����             - < _ %          z  n
       $       ���       ���� � �������������          ����             0 ? d '          �  "       $       ���       ���� � �������������          ����             3 B i )          �  �       $       ���       ���� � �������������          ����             6 E n +           .  �       $       ���       ���� � �������������          ����             9 H s -       !   j  >       $	       ���       ���� � �������������         ����             & 4 `        6   Z  h       %        ���        ���� � �������������         ����  	 
          ) 8 e        :   �  �       %       ���        ���� � �������������         ����             , < j        >     8       %       ���        ���� � �������������         ����             / @ o "       A   h  �       %       ���       ���� � �������������         ����             2 D t %       E   �         %       ���       ���� � �������������         ����             5 H y (       H     p       %       ���       ���� � �������������         ����             8 L ~ +       L   v  �       %       ���       ���� � �������������         ����             ; P � .       P   �  @       %       ���       ���� � �������������         ����             > T � 1       S   *  �        %       ���       ���� � �������������         ����             A X � 4       W   �  "       %	       ���       ���� � �������������         ����  
           . E y !          �	  �1       &        ���        ���� � �������������         ����             1 I  $       �   d
  �3       &       ���        ���� � �������������         ����             4 M � '       �   �
  L6       &       ���        ���� � �������������         ����             7 Q � *       �   T  �8       &       ���       ���� � �������������         ����             : U � -       �   �  �:       &       ���       ���� � �������������         ����             = Y � 0       �   D  T=       &       ���       ���� � �������������         ����             @ ] � 3       �   �  �?       &       ���       ���� � �������������         ����             C a � 6       �   4  B       &       ���       ���� � �������������         ����             F e � 9       �   �  \D       &       ���       ���� � �������������         ����             I i � <       �   $  �F       &	       ���       ���� � �������������         ����             5 U � (       �     `       '        ���        ���� � �������������         ����             8 Y � +       �   �  �c       '       ���        ���� � �������������         ����             ; ] � .         0   g       '       ���        ���� � �������������         ����             > a � 1         �  �j       '       ���       ���� � �������������         ����             A e � 4         \  (n       '       ���       ���� � �������������         ����             D i � 7       #  �  �q       '       ���       ���� � �������������         ����             G m � :       ,  �  0u       '       ���       ���� � �������������         ����             J q � =       5    �x       '       ���       ���� � �������������         ����             M u � @       >  �  8|    
   '       ���       ���� � �������������         ����              P y � C       G  J  �    	   '	       ���       ���� � �������������          ����             
  %        !   �  /       �        ���        ���� � �������������          ����               *        (   �  �       �       ���        ���� � �������������          ����               /        )            �       ���        ���� � �������������          ����                4        )   *  T       �       ���       ���� � �������������          ����  	 
           # 9        *   H  �       �       ���       ���� � �������������          ����              & >        +   f  �       �       ���       ���� � �������������          ����              ) C        +   �         �       ���       ���� � �������������          ����              , H        ,   �  D       �       ���       ���� � �������������          ����              / M         ,   �  �       �       ���       ���� � �������������          ����              2 R "       -   �  �       �	       ���       ���� � �������������          ����             	  @        G   V	         �        ���        ���� � �������������          ����              " E        I   �	  �       �       ���        ���� � �������������          ����   	           % J        K   �	  j       �       ���        ���� � �������������          ����  
            ( O        M   

         �       ���       ���� � �������������          ����              + T        N   F
  �       �       ���       ���� � �������������          ����              . Y        P   �
  �       �       ���       ���� � �������������          ����              1 ^        R   �
  :        �       ���       ���� � �������������          ����              4 c        T   �
  �        �       ���       ���� � �������������          ����             ! 7 h        V   6  �!       �       ���       ���� � �������������          ����             $ : m !       W   r  V"       �	       ���       ���� � �������������          ����              & Z        ~   b  �1       �        ���        ���� � �������������         ����  	 
           * _        �   �  �2       �       ���        ���� � �������������         ����              . d        �     X4       �       ���        ���� � �������������         ����              2 i        �   p  �5       �       ���       ���� � �������������         ����              6 n        �   �  (7       �       ���       ���� � �������������         ����               : s        �   $  �8       �       ���       ���� � �������������         ����             # > x        �   ~  �9       �       ���       ���� � �������������         ����             & B } "       �   �  `;       �       ���       ���� � �������������         ����             ) F � %       �   2  �<       �       ���       ���� � �������������         ����             , J � (       �   �  0>       �	       ���       ���� � �������������          ����  
            7 s        �   �  �T       �        ���        ���� � �������������         ����              ; y        �   l  W       �       ���        ���� � �������������         ����              ?         �   �  tY       �       ���        ���� � �������������         ����             " C �        �   \  �[       �       ���       ���� � �������������         ����             % G � !       �   �  $^       �       ���       ���� � �������������         ����             ( K � $       �   L  |`       �       ���       ���� � �������������         ����             + O � '       �   �  �b       �       ���       ���� � �������������         ����             . S � *         <  ,e       �       ���       ���� � �������������         ����             1 W � -       	  �  �g       �       ���       ���� � �������������         ����             4 [ � 0         ,  �i       �	       ���       ���� � �������������          ����               G �        b    H�       �        ���        ���� � �������������         ����             # K �        k  �  ̍       �       ���        ���� � �������������         ����             & O � "       t  8  P�       �       ���        ���� � �������������         ����             ) S � %       }  �  Ԕ       �       ���       ���� � �������������         ����             , W � (       �  d  X�       �       ���       ���� � �������������         ����             / [ � +       �  �  ܛ       �       ���       ���� � �������������         ����             2 _ � .       �  �  `�       �       ���       ���� � �������������         ����             5 c � 1       �  &  �       �       ���       ���� � �������������         ����             8 g � 4       �  �  h�    
   �       ���       ���� � �������������         ����              ; k � 7       �  R  �    	   �	       ���       ���� � �������������          ����             % 2 @ +          @  �       �         ���        ���� � �������������          ����             ' 5 E -           ^  �       �        ���        ���� � �������������          ����             ) 8 J /       !   |  �       �        ���        ���� � �������������          ����   	          + ; O 1       !   �  4       �        ���       ���� � �������������          ����  
           - > T 3       "   �  p       �        ���       ���� � �������������          ����             / A Y 5       #   �  �       �        ���       ���� � �������������          ����             1 D ^ 7       #   �  �       �        ���       ���� � �������������          ����             3 G c 9       $     $       �        ���       ���� � �������������          ����             5 J h ;       $   0  `       �        ���       ���� � �������������          ����             7 M m =       %   N  �       �	        ���       ���� � �������������          ����             $ : [ *       ;   �  R       �        ���        ���� � �������������          ����             ' = ` ,       =            �       ���        ���� � �������������          ����  	 
          * @ e .       ?   >  �       �       ���        ���� � �������������          ����             - C j 0       A   z  n       �       ���       ���� � �������������          ����             0 F o 2       B   �  "       �       ���       ���� � �������������          ����             3 I t 4       D   �  �       �       ���       ���� � �������������          ����             6 L y 6       F   .	  �       �       ���       ���� � �������������          ����             9 O ~ 8       H   j	  >       �       ���       ���� � �������������          ����             < R � :       J   �	  �       �       ���       ���� � �������������          ����             ? U � <       K   �	  �       �	       ���       ���� � �������������         ����   	          , A u (       n   �
  H+       �        ���        ���� � �������������         ����  
           / E z +       r   ,  �,       �       ���        ���� � �������������         ����             2 I  .       v   �  .       �       ���        ���� � �������������         ����             5 M � 1       y   �  �/       �       ���       ���� � �������������         ����             8 Q � 4       }   :  �0       �       ���       ���� � �������������         ����             ; U � 7       �   �  P2       �       ���       ���� � �������������         ����             > Y � :       �   �  �3       �       ���       ���� � �������������         ����             A ] � =       �   H   5       �       ���       ���� � �������������         ����             D a � @       �   �  �6       �       ���       ���� � �������������         ����             G e � C       �   �  �7       �	       ���       ���� � �������������         ����             4 R � 0       �   d  �L       �        ���        ���� � �������������         ����             7 V � 3       �   �  LO       �       ���        ���� � �������������         ����             : Z � 6       �   T  �Q       �       ���        ���� � �������������         ����             = ^ � 9       �   �  �S       �       ���       ���� � �������������         ����             @ b � <       �   D  TV       �       ���       ���� � �������������         ����             C f � ?       �   �  �X       �       ���       ���� � �������������         ����             F j � B       �   4  [       �       ���       ���� � �������������         ����             I n � E       �   �  \]       �       ���       ���� � �������������         ����             L r � H       �   $  �_       �       ���       ���� � �������������         ����             O v � K       �   �  b       �	       ���       ���� � �������������         ����             ; b � 7       J  |  �       �        ���        ���� � �������������         ����             > f � :       S    l�       �       ���        ���� � �������������         ����             A j � =       \  �  ��       �       ���        ���� � �������������         ����             D n � @       e  >  t�       �       ���       ���� � �������������         ����             G r � C       n  �  ��       �       ���       ���� � �������������         ����             J v � F       w  j  |�       �       ���       ���� � �������������         ����             M z � I       �      �       �       ���       ���� � �������������         ����             P ~ � L       �  �  ��       �       ���       ���� � �������������         ����             S � � O       �  ,  �    
   �       ���       ���� � �������������         ����    !          V � � R       �  �  ��    	   �	       ���       ���� � �������������          ����              ) 7 "          �  F       U        ���        ���� � �������������          ����              , < $          �  �	       U       ���        ���� � �������������          ����               / A &          �  �	       U       ���        ���� � �������������          ����             " 2 F (          
  
       U       ���       ���� � �������������          ����  	 
          $ 5 K *          (  P
       U       ���       ���� � �������������          ����             & 8 P ,          F  �
       U       ���       ���� � �������������          ����             ( ; U .          d  �
       U       ���       ���� � �������������          ����             * > Z 0          �         U       ���       ���� � �������������          ����             , A _ 2          �  @       U       ���       ���� � �������������          ����             . D d 4          �  |       U	       ���       ���� � �������������          ����              1 R !       /   6  �       V        ���        ���� � �������������          ����              4 W #       1   r  V       V       ���        ���� � �������������          ����   	          ! 7 \ %       3   �  
       V       ���        ���� � �������������          ����  
           $ : a '       5   �  �       V       ���       ���� � �������������          ����             ' = f )       6   &  r       V       ���       ���� � �������������          ����             * @ k +       8   b  &       V       ���       ���� � �������������          ����             - C p -       :   �  �       V       ���       ���� � �������������          ����             0 F u /       <   �  �       V       ���       ���� � �������������          ����             3 I z 1       >     B       V       ���       ���� � �������������          ����             6 L  3       ?   R  �       V	       ���       ���� � �������������          ����             # 8 l        ^   B	  %       W        ���        ���� � �������������         ����  	 
          & < q "       b   �	  p&       W       ���        ���� � �������������         ����             ) @ v %       f   �	  �'       W       ���        ���� � �������������         ����             , D { (       i   P
  @)       W       ���       ���� � �������������         ����             / H � +       m   �
  �*       W       ���       ���� � �������������         ����             2 L � .       p     ,       W       ���       ���� � �������������         ����             5 P � 1       t   ^  x-       W       ���       ���� � �������������         ����             8 T � 4       x   �  �.       W       ���       ���� � �������������         ����             ; X � 7       {     H0       W       ���       ���� � �������������         ����             > \ � :          l  �1       W	       ���       ���� � �������������          ����  
           + I � '       �   �  $E       X        ���        ���� � �������������         ����             . M � *       �   L  |G       X       ���        ���� � �������������         ����             1 Q � -       �   �  �I       X       ���        ���� � �������������         ����             4 U � 0       �   <  ,L       X       ���       ���� � �������������         ����             7 Y � 3       �   �  �N       X       ���       ���� � �������������         ����             : ] � 6       �   ,  �P       X       ���       ���� � �������������         ����             = a � 9       �   �  4S       X       ���       ���� � �������������         ����             @ e � <       �     �U       X       ���       ���� � �������������         ����             C i � ?       �   �  �W       X       ���       ���� � �������������         ����             F m � B       �     <Z       X	       ���       ���� � �������������          ����             2 Y � .       2  �  �w       Y        ���        ���� � �������������         ����             5 ] � 1       ;  �  {       Y       ���        ���� � �������������         ����             8 a � 4       D    �~       Y       ���        ���� � �������������         ����             ; e � 7       M  �  �       Y       ���       ���� � �������������         ����             > i � :       V  D  ��       Y       ���       ���� � �������������         ����             A m � =       _  �  �       Y       ���       ���� � �������������         ����             D q � @       h  p  ��       Y       ���       ���� � �������������         ����             G u � C       q    $�       Y       ���       ���� � �������������         ����             J y � F       z  �  ��    
   Y       ���       ���� � �������������         ����              M } � I       �  2  ,�    	   Y	       ���       ���� � �������������          H g                    
       �����   �        
      ��' ���        ����   ����������������        I g                          ����B  �              ��' ���        ����   ����������������        J g                  $        ����[  l              ��' ���        ����   ����������������        K g                " & 9        ����'  �#              ��' ���        ����   ����������������        L g                2 6 P !       �����
  �?              ��' ���        ����   ����������������        M g                A H i (       �����  �g              ��' ���        ����   ����������������         g                Q W  1       �����  �              ��' ���        ����   ����������������         g                c d � :       ����U  ��              ��' ���        ����   ����������������        N g                k l � B       �����  @<             ��' ���        ����	   ����������������        O g                { } � I       �����&  ʨ             ��' ���        ����
   ����������������        P g                � � � T       ����O.  �+             ��' ���        ����   ����������������        Q g                � � � ^       �����6  �             ��' ���        ����   ����������������        R g                � � k       �����?  }             ��' ���        ����   ����������������        S g                � � &~       �����I  �O             ��' ���        ����   ����������������        T g                � � I�       ����T  A             ��' ���        ����   ����������������        U g                � q�       ����A_  QS             ��' ���        ����   ����������������        V g                �  ��       ����$k  ��             ��' ���        ����   ����������������        W g                A��       �����w  ��             ��' ���        ����   ����������������        X g                 d�       �����  <d
             ��' ���        ����   ����������������        Y g                9�C�       ������  �             ��' ���        ����   ����������������        Z g                R��      ������  ��             ��' ���        ����   ����������������        [ g                j��      �����  p�             ��' ���        ����   ����������������        \ g                ���.      ����%�  x              ��' ���        ����   ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ���        ������  ����������������       ����� ��                            ����'   N        �      ��R ��         ������  ����������������       ����   2 3          Z� h \       �  �G  z   	         
  ��        ����
 � �����  �  �         ����   4 5          a� l `         �H  ^!           
  ��        ����
 � �����  �  �         ����   6 7          h� p d       $  J  B.           
  ��        ����
 � �����  �  �         ����   9 :          o� t h       E  2K  &;           
  ��       ����
 � �����  �  �         ����   ; <          v� x l       f  ^L  
H           
  ��       ����
 � �����  �  �         ����   = >          }� | p       �  �M  �T           
  ��       ����
 � �����  �  �         ����   ? @          �� � t       �  �N  �a           
  ��       ����
 � �����  �  �         ����   A B          �� � x       �  �O  �n   ��       
  ��       ����
 � �����  �  �         ����   D E          �� � |       �  Q  �{   ��       
  ��       ����
 � �����  �  �         ����   F G          �� � �       	  :R  ~�   ��  	     
  ��       ����
 7  �  �  �         ����   < =          � d           	      �        %        ��        ����c   �������������         ����   > ?          � g              >  |        %       ��        ����c   �������������         ����   @ A          � j              \  �        %       ��        ����c   �������������         ����   B C          � m              z  �        %       ��       ����c   �������������         ����   D E          � p              �  0        %       ��       ����c   �������������         ����   F G          � s              �  l        %       ��       ����c   �������������         ����   H I          � v              �  �        %       ��       ����c   �������������         ����   J K          � y              �  �        %       ��       ����c   �������������         ����   L M          � |                         %       ��       ����c   �������������         ����   N O          �               .  \        %	       ��       ����c   �������������         ����   ' (          � � Sb       �  �G  z   	   3      
  ��        ����
 � �����  �  �         ����   ) *          � � Zf         �H  ^!      3     
  ��        ����
 � �����  �  �         ����   + ,          � � aj       $  J  B.      3     
  ��        ����
 � �����  �  �         ����   - .          � � hn       E  2K  &;      3     
  ��       ����
 � �����  �  �         ����   / 0          � � or       f  ^L  
H      3     
  ��       ����
 � �����  �  �         ����   1 2          � � vv       �  �M  �T      3     
  ��       ����
 � �����  �  �         ����   4 5          � � }z       �  �N  �a      3     
  ��       ����
 � �����  �  �         ����   6 7          � � �~       �  �O  �n   ��  3     
  ��       ����
 � �����  �  �         ����   8 9          � � ��       �  Q  �{   ��  3     
  ��       ����
 � �����  �  �         ����   : ;          � � ��       	  :R  ~�   ��  3	     
  ��       ����
 7  �  �  �         ����   2 3            d �         	      �        9        ��        ����c   �������������         ����   4 5            g �            >  |        9       ��        ����c   �������������         ����   6 7            j �            \  �        9       ��        ����c   �������������         ����   8 9            m �            z  �        9       ��       ����c   �������������         ����   : ;            p �            �  0        9       ��       ����c   �������������         ����   < =            s �            �  l        9       ��       ����c   �������������         ����   > ?            v �            �  �        9       ��       ����c   �������������         ����   @ A            y �            �  �        9       ��       ����c   �������������         ����   B C            | �                       9       ��       ����c   �������������         ����   D E             �            .  \        9	       ��       ����c   �������������         ����   & '          [ ]       �  �G  z   	   G      
  ��        ����
 � �����  �  �         ����   ( )          _ a         �H  ^!      G     
  ��        ����
 � �����  �  �         ����   * +          "c "e       $  J  B.      G     
  ��        ����
 � �����  �  �         ����   , -          (g (i       E  2K  &;      G     
  ��       ����
 � �����  �  �         ����   . /          .k .m       f  ^L  
H      G     
  ��       ����
 � �����  �  �         ����   0 1          4o 4q       �  �M  �T      G     
  ��       ����
 � �����  �  �         ����   3 4          :s :u       �  �N  �a      G     
  ��       ����
 � �����  �  �         ����   5 6          @w @y       �  �O  �n   ��  G     
  ��       ����
 � �����  �  �         ����   7 8          F{ F}       �  Q  �{   ��  G     
  ��       ����
 � �����  �  �         ����   9 :          L L�       	  :R  ~�   ��  G	     
  ��       ����
 7  �  �  �         ����   1 2          �   �         	      �        M        ��        ����c   �������������         ����   3 4          �   �            >  |        M       ��        ����c   �������������         ����   5 6          �   �            \  �        M       ��        ����c   �������������         ����   7 8          �   �            z  �        M       ��       ����c   �������������         ����   9 :          �   �            �  0        M       ��       ����c   �������������         ����   ; <          �   �            �  l        M       ��       ����c   �������������         ����   = >          �   �            �  �        M       ��       ����c   �������������         ����   ? @          �   �            �  �        M       ��       ����c   �������������         ����   A B          �   �                       M       ��       ����c   �������������         ����   C D          �   �            .  \        M	       ��       ����c   �������������         ����  0 1          E� h \       �  �E  ��   	   �      
  ��        ����
 � �����  �  �         ����  2 3          L� l `       �  �F  �      �     
  ��        ����
 � �����  �  �         ����  4 5          S� p d       �  H  �      �     
  ��        ����
 � �����  �  �         ����  7 8          Z� t h         >I  �%      �     
  ��       ����
 � �����  �  �         ����  9 :          a� x l       /  jJ  �2      �     
  ��       ����
 � �����  �  �         ����  ; <          h� | p       P  �K  r?      �     
  ��       ����
 � �����  �  �         ����  = >          o� � t       q  �L  VL      �     
  ��       ����
 � �����  �  �         ����  ? @          v� � x       �  �M  :Y   ��  �     
  ��       ����
 � �����  �  �         ����  B C          }� � |       �  O  f   ��  �     
  ��       ����
 � �����  �  �         ����  D E          �� � �       �  FP  s   ��  �	     
  ��       ����
 7  �  �  �         ����  : ;          � d              ,  h        �        ��        ����c   �������������         ����  < =          � g              J  �        �       ��        ����c   �������������         ����  > ?          � j              h  �        �       ��        ����c   �������������         ����  @ A          � m              �          �       ��       ����c   �������������         ����  B C          � p              �  H        �       ��       ����c   �������������         ����  D E          � s           	   �  �        �       ��       ����c   �������������         ����  F G          � v           	   �  �        �       ��       ����c   �������������         ����  H I          � y           
   �  �        �       ��       ����c   �������������         ����  J K          � |           
     8        �       ��       ����c   �������������         ����  L M          �               :  t        �	       ��       ����c   �������������         ����  & '          q � >b       �  �E  ��   	   �      
  ��	        ����
 � �����  �  �         ����  ( )          v � Ef       �  �F  �      �     
  ��	        ����
 � �����  �  �         ����  * +          { � Lj       �  H  �      �     
  ��	        ����
 � �����  �  �         ����  , -          � � Sn         >I  �%      �     
  ��	       ����
 � �����  �  �         ����  . /          � � Zr       /  jJ  �2      �     
  ��	       ����
 � �����  �  �         ����  0 1          � � av       P  �K  r?      �     
  ��	       ����
 � �����  �  �         ����  3 4          � � hz       q  �L  VL      �     
  ��	       ����
 � �����  �  �         ����  5 6          � � o~       �  �M  :Y   ��  �     
  ��	       ����
 � �����  �  �         ����  7 8          � � v�       �  O  f   ��  �     
  ��	       ����
 � �����  �  �         ����  9 :          � � }�       �  FP  s   ��  �	     
  ��	       ����
 7  �  �  �         ����  1 2            d �            ,  h        �        ��
        ����c   �������������         ����  3 4            g �            J  �        �       ��
        ����c   �������������         ����  5 6            j �            h  �        �       ��
        ����c   �������������         ����  7 8            m �            �          �       ��
       ����c   �������������         ����  9 :            p �            �  H        �       ��
       ����c   �������������         ����  ; <            s �         	   �  �        �       ��
       ����c   �������������         ����  = >            v �         	   �  �        �       ��
       ����c   �������������         ����  ? @            y �         
   �  �        �       ��
       ����c   �������������         ����  A B            | �         
     8        �       ��
       ����c   �������������         ����  C D             �            :  t        �	       ��
       ����c   �������������         ����  % &          [ ]       �  �E  ��   	   �      
  ��        ����
 � �����  �  �         ����  ' (          _ a       �  �F  �      �     
  ��        ����
 � �����  �  �         ����  ) *          c e       �  H  �      �     
  ��        ����
 � �����  �  �         ����  + ,          g i         >I  �%      �     
  ��       ����
 � �����  �  �         ����  - .          k m       /  jJ  �2      �     
  ��       ����
 � �����  �  �         ����  / 0          o q       P  �K  r?      �     
  ��       ����
 � �����  �  �         ����  2 3          %s %u       q  �L  VL      �     
  ��       ����
 � �����  �  �         ����  4 5          +w +y       �  �M  :Y   ��  �     
  ��       ����
 � �����  �  �         ����  6 7          1{ 1}       �  O  f   ��  �     
  ��       ����
 � �����  �  �         ����  8 9          7 7�       �  FP  s   ��  �	     
  ��       ����
 7  �  �  �         ����  0 1          �   �            ,  h        �        ��        ����c   �������������         ����  2 3          �   �            J  �        �       ��        ����c   �������������         ����  4 5          �   �            h  �        �       ��        ����c   �������������         ����  6 7          �   �            �          �       ��       ����c   �������������         ����  8 9          �   �            �  H        �       ��       ����c   �������������         ����  : ;          �   �         	   �  �        �       ��       ����c   �������������         ����  < =          �   �         	   �  �        �       ��       ����c   �������������         ����  > ?          �   �         
   �  �        �       ��       ����c   �������������         ����  @ A          �   �         
     8        �       ��       ����c   �������������         ����  B C          �   �            :  t        �	       ��       ����c   �������������         ����  1 2          R� h \       �  VE  ��   	   �      
  ��        ����
 � �����  �  �         ����  3 4          Y� l `       �  �F  �      �     
  ��        ����
 � �����  �  �         ����  5 6          `� p d       �  �G  z      �     
  ��        ����
 � �����  �  �         ����  8 9          g� t h         �H  ^!      �     
  ��       ����
 � �����  �  �         ����  : ;          n� x l       $  J  B.      �     
  ��       ����
 � �����  �  �         ����  < =          u� | p       E  2K  &;      �     
  ��       ����
 � �����  �  �         ����  > ?          |� � t       f  ^L  
H      �     
  ��       ����
 � �����  �  �         ����  @ A          �� � x       �  �M  �T   ��  �     
  ��       ����
 � �����  �  �         ����  C D          �� � |       �  �N  �a   ��  �     
  ��       ����
 � �����  �  �         ����  E F          �� � �       �  �O  �n   ��  �	     
  ��       ����
 7  �  �  �         ����  ; <          � d              �   �         �        ��        ����c   �������������         ����  = >          � g              �   �        �       ��        ����c   �������������         ����  ? @          � j                        �       ��        ����c   �������������         ����  A B          � m              "  D        �       ��       ����c   �������������         ����  C D          � p              @  �        �       ��       ����c   �������������         ����  E F          � s              ^  �        �       ��       ����c   �������������         ����  G H          � v              |  �        �       ��       ����c   �������������         ����  I J          � y              �  4        �       ��       ����c   �������������         ����  K L          � |              �  p        �       ��       ����c   �������������         ����  M N          �            	   �  �        �	       ��       ����c   �������������         ����  & '          ~ � Kb       �  VE  ��   	   
      
  ��        ����
 � �����  �  �         ����  ( )          � � Rf       �  �F  �      
     
  ��        ����
 � �����  �  �         ����  * +          � � Yj       �  �G  z      
     
  ��        ����
 � �����  �  �         ����  , -          � � `n         �H  ^!      
     
  ��       ����
 � �����  �  �         ����  . /          � � gr       $  J  B.      
     
  ��       ����
 � �����  �  �         ����  0 1          � � nv       E  2K  &;      
     
  ��       ����
 � �����  �  �         ����  3 4          � � uz       f  ^L  
H      
     
  ��       ����
 � �����  �  �         ����  5 6          � � |~       �  �M  �T   ��  
     
  ��       ����
 � �����  �  �         ����  7 8          � � ��       �  �N  �a   ��  
     
  ��       ����
 � �����  �  �         ����  9 :          � � ��       �  �O  �n   ��  
	     
  ��       ����
 7  �  �  �         ����  1 2            d �            �   �                 ��        ����c   �������������         ����  3 4            g �            �   �               ��        ����c   �������������         ����  5 6            j �                             ��        ����c   �������������         ����  7 8            m �            "  D               ��       ����c   �������������         ����  9 :            p �            @  �               ��       ����c   �������������         ����  ; <            s �            ^  �               ��       ����c   �������������         ����  = >            v �            |  �               ��       ����c   �������������         ����  ? @            y �            �  4               ��       ����c   �������������         ����  A B            | �            �  p               ��       ����c   �������������         ����  C D             �         	   �  �        	       ��       ����c   �������������         ����  % &          [ ]       �  VE  ��   	         
  ��        ����
 � �����  �  �         ����  ' (          _ a       �  �F  �           
  ��        ����
 � �����  �  �         ����  ) *          c e       �  �G  z           
  ��        ����
 � �����  �  �         ����  + ,           g  i         �H  ^!           
  ��       ����
 � �����  �  �         ����  - .          &k &m       $  J  B.           
  ��       ����
 � �����  �  �         ����  / 0          ,o ,q       E  2K  &;           
  ��       ����
 � �����  �  �         ����  2 3          2s 2u       f  ^L  
H           
  ��       ����
 � �����  �  �         ����  4 5          8w 8y       �  �M  �T   ��       
  ��       ����
 � �����  �  �         ����  6 7          >{ >}       �  �N  �a   ��       
  ��       ����
 � �����  �  �         ����  8 9          D D�       �  �O  �n   ��  	     
  ��       ����
 7  �  �  �         ����  0 1          �   �            �   �         !        ��        ����c   �������������         ����  2 3          �   �            �   �        !       ��        ����c   �������������         ����  4 5          �   �                      !       ��        ����c   �������������         ����  6 7          �   �            "  D        !       ��       ����c   �������������         ����  8 9          �   �            @  �        !       ��       ����c   �������������         ����  : ;          �   �            ^  �        !       ��       ����c   �������������         ����  < =          �   �            |  �        !       ��       ����c   �������������         ����  > ?          �   �            �  4        !       ��       ����c   �������������         ����  @ A          �   �            �  p        !       ��       ����c   �������������         ����  B C          �   �         	   �  �        !	       ��       ����c   �������������         ����  0 1          @� h \       f  ^L  
H   	   _      
  ��        ����
 � �����  �  �         ����  2 3          G� l `       �  �M  �T      _     
  ��        ����
 � �����  �  �         ����  4 5          N� p d       �  �N  �a      _     
  ��        ����
 � �����  �  �         ����  7 8          U� t h       �  �O  �n      _     
  ��       ����
 � �����  �  �         ����  9 :          \� x l       �  Q  �{      _     
  ��       ����
 � �����  �  �         ����  ; <          c� | p       	  :R  ~�      _     
  ��       ����
 � �����  �  �         ����  = >          j� � t       ,	  fS  b�      _     
  ��       ����
 � �����  �  �         ����  ? @          q� � x       M	  �T  F�   ��  _     
  ��       ����
 � �����  �  �         ����  B C          x� � |       n	  �U  *�   ��  _     
  ��       ����
 � �����  �  �         ����  D E          � � �       �	  �V  �   ��  _	     
  ��       ����
 7  �  �  �         ����  : ;          � d           !   �  /        e        ��        ����c   �������������         ����  < =          � g           (   �  �        e       ��        ����c   �������������         ����  > ?          � j           )             e       ��        ����c   �������������         ����  @ A          � m           )   *  T        e       ��       ����c   �������������         ����  B C          � p           *   H  �        e       ��       ����c   �������������         ����  D E          � s           +   f  �        e       ��       ����c   �������������         ����  F G          � v           +   �          e       ��       ����c   �������������         ����  H I          � y           ,   �  D        e       ��       ����c   �������������         ����  J K          � |           ,   �  �        e       ��       ����c   �������������         ����  L M          �            -   �  �        e	       ��       ����c   �������������         ����  & '          l � 9b       f  ^L  
H   	   p      
  ��        ����
 � �����  �            ����  ( )          q � @f       �  �M  �T      p     
  ��        ����
 � �����  �            ����  * +          v � Gj       �  �N  �a      p     
  ��        ����
 � �����  �            ����  , -          { � Nn       �  �O  �n      p     
  ��       ����
 � �����  �            ����  . /          � � Ur       �  Q  �{      p     
  ��       ����
 � �����  �            ����  0 1          � � \v       	  :R  ~�      p     
  ��       ����
 � �����  �            ����  3 4          � � cz       ,	  fS  b�      p     
  ��       ����
 � �����  �            ����  5 6          � � j~       M	  �T  F�   ��  p     
  ��       ����
 � �����  �            ����  7 8          � � q�       n	  �U  *�   ��  p     
  ��       ����
 � �����  �            ����  9 :          � � x�       �	  �V  �   ��  p	     
  ��       ����
 7  �  �            ����  1 2            d �         !   �  /        v        ��        ����c   ������������         ����  3 4            g �         (   �  �        v       ��        ����c   ������������         ����  5 6            j �         )             v       ��        ����c   ������������         ����  7 8            m �         )   *  T        v       ��       ����c   ������������         ����  9 :            p �         *   H  �        v       ��       ����c   ������������         ����  ; <            s �         +   f  �        v       ��       ����c   ������������         ����  = >            v �         +   �          v       ��       ����c   ������������         ����  ? @            y �         ,   �  D        v       ��       ����c   ������������         ����  A B            | �         ,   �  �        v       ��       ����c   ������������         ����  C D             �         -   �  �        v	       ��       ����c   ������������         ����  % &          � [ � ]       f  ^L  
H   	   �      
  ��        ����
 � �����  �           ����  ' (          _ a       �  �M  �T      �     
  ��        ����
 � �����  �           ����  ) *          c e       �  �N  �a      �     
  ��        ����
 � �����  �           ����  + ,          g i       �  �O  �n      �     
  ��       ����
 � �����  �           ����  - .          k m       �  Q  �{      �     
  ��       ����
 � �����  �           ����  / 0          o q       	  :R  ~�      �     
  ��       ����
 � �����  �           ����  2 3           s  u       ,	  fS  b�      �     
  ��       ����
 � �����  �           ����  4 5          &w &y       M	  �T  F�   ��  �     
  ��       ����
 � �����  �           ����  6 7          ,{ ,}       n	  �U  *�   ��  �     
  ��       ����
 � �����  �           ����  8 9          2 2�       �	  �V  �   ��  �	     
  ��       ����
 7  �  �           ����  1 2          �   �         !   �  /        �        ��        ����c   ������������         ����  3 4          �   �         (   �  �        �       ��        ����c   ������������         ����  5 6          �   �         )             �       ��        ����c   ������������         ����  7 8          �   �         )   *  T        �       ��       ����c   ������������         ����  9 :          �   �         *   H  �        �       ��       ����c   ������������         ����  ; <          �   �         +   f  �        �       ��       ����c   ������������         ����  = >          �   �         +   �          �       ��       ����c   ������������         ����  ? @          �   �         ,   �  D        �       ��       ����c   ������������         ����  A B          �   �         ,   �  �        �       ��       ����c   ������������         ����  C D          �   �         -   �  �        �	       ��       ����c   ������������         ����  3 4          g� h \       :  �J  �6   	   �      	  ��        ����
 � �����  �           ����  5 6          n� l `       [  �K  �C      �     	  ��        ����
 � �����  �           ����  7 8          u� p d       |  &M  �P      �     	  ��        ����
 � �����  �           ����  : ;          |� t h       �  RN  �]      �     	  ��       ����
 � �����  �           ����  < =          �� x l       �  ~O  jj      �     	  ��       ����
 � �����  �           ����  > ?          �� | p       �  �P  Nw      �     	  ��       ����
 � �����  �           ����  @ A          �� � t        	  �Q  2�      �     	  ��       ����
 � �����  �           ����  B C          �� � x       !	  S  �   ��  �     	  ��       ����
 � �����  �           ����  E F          �� � |       B	  .T  ��   ��  �     	  ��       ����
 � �����  �           ����  G H          �� � �       c	  ZU  ު   ��  �	     	  ��       ����
 7  �  �           ����  = >          � d              @  �        �        ��        ����c   ������������         ����  ? @          � g               ^  �        �       ��        ����c   ������������         ����  A B          � j           !   |  �        �       ��        ����c   ������������         ����  C D          � m           !   �  4        �       ��       ����c   ������������         ����  E F          � p           "   �  p        �       ��       ����c   ������������         ����  G H          � s           #   �  �        �       ��       ����c   ������������         ����  I J          � v           #   �  �        �       ��       ����c   ������������         ����  K L          � y           $     $        �       ��       ����c   ������������         ����  M N          � |           $   0  `        �       ��       ����c   ������������         ����  O P          �            %   N  �        �	       ��       ����c   ������������         ����  ' (          � � `b       :  �J  �6   	   �      	  ��        ����
 � �����  �           ����  ) *          � � gf       [  �K  �C      �     	  ��        ����
 � �����  �           ����  + ,          � � nj       |  &M  �P      �     	  ��        ����
 � �����  �           ����  - .          � � un       �  RN  �]      �     	  ��       ����
 � �����  �           ����  / 0          � � |r       �  ~O  jj      �     	  ��       ����
 � �����  �           ����  1 2          � � �v       �  �P  Nw      �     	  ��       ����
 � �����  �           ����  4 5          � � �z        	  �Q  2�      �     	  ��       ����
 � �����  �           ����  6 7          � � �~       !	  S  �   ��  �     	  ��       ����
 � �����  �           ����  8 9          � � ��       B	  .T  ��   ��  �     	  ��       ����
 � �����  �           ����  : ;          � � ��       c	  ZU  ު   ��  �	     	  ��       ����
 7  �  �           ����  2 3            d �            @  �        �        ��        ����c   ������������         ����  4 5            g �             ^  �        �       ��        ����c   ������������         ����  6 7            j �         !   |  �        �       ��        ����c   ������������         ����  8 9            m �         !   �  4        �       ��       ����c   ������������         ����  : ;            p �         "   �  p        �       ��       ����c   ������������         ����  < =            s �         #   �  �        �       ��       ����c   ������������         ����  > ?            v �         #   �  �        �       ��       ����c   ������������         ����  @ A            y �         $     $        �       ��       ����c   ������������         ����  B C            | �         $   0  `        �       ��       ����c   ������������         ����  D E             �         %   N  �        �	       ��       ����c   ������������         ����  & '          #[ #]       :  �J  �6   	   �      	  ��        ����
 � �����  �           ����  ( )          )_ )a       [  �K  �C      �     	  ��        ����
 � �����  �           ����  * +          /c /e       |  &M  �P      �     	  ��        ����
 � �����  �           ����  , -          5g 5i       �  RN  �]      �     	  ��       ����
 � �����  �           ����  . /          ;k ;m       �  ~O  jj      �     	  ��       ����
 � �����  �           ����  0 1          Ao Aq       �  �P  Nw      �     	  ��       ����
 � �����  �           ����  3 4          Gs Gu        	  �Q  2�      �     	  ��       ����
 � �����  �           ����  5 6          Mw My       !	  S  �   ��  �     	  ��       ����
 � �����  �           ����  7 8          S{ S}       B	  .T  ��   ��  �     	  ��       ����
 � �����  �           ����  9 :          Y Y�       c	  ZU  ު   ��  �	     	  ��       ����
 7  �  �           ����  1 2          �   �            @  �        �        ��        ����c   ������������	         ����  3 4          �   �             ^  �        �       ��        ����c   ������������	         ����  5 6          �   �         !   |  �        �       ��        ����c   ������������	         ����  7 8          �   �         !   �  4        �       ��       ����c   ������������	         ����  9 :          �   �         "   �  p        �       ��       ����c   ������������	         ����  ; <          �   �         #   �  �        �       ��       ����c   ������������	         ����  = >          �   �         #   �  �        �       ��       ����c   ������������	         ����  ? @          �   �         $     $        �       ��       ����c   ������������	         ����  A B          �   �         $   0  `        �       ��       ����c   ������������	         ����  C D          �   �         %   N  �        �	       ��       ����c   ������������	         ����  1 2          M� h \         >I  �%   	   +      
  ��        ����
 � �����  �  
         ����  3 4          T� l `       /  jJ  �2      +     
  ��        ����
 � �����  �  
         ����  5 6          [� p d       P  �K  r?      +     
  ��        ����
 � �����  �  
         ����  8 9          b� t h       q  �L  VL      +     
  ��       ����
 � �����  �  
         ����  : ;          i� x l       �  �M  :Y      +     
  ��       ����
 � �����  �  
         ����  < =          p� | p       �  O  f      +     
  ��       ����
 � �����  �  
         ����  > ?          w� � t       �  FP  s      +     
  ��       ����
 � �����  �  
         ����  @ A          ~� � x       �  rQ  �   ��  +     
  ��       ����
 � �����  �  
         ����  C D          �� � |       	  �R  ʌ   ��  +     
  ��       ����
 � �����  �  
         ����  E F          �� � �       7	  �S  ��   ��  +	     
  ��       ����
 7  �  �  
         ����  ; <          � d              �  F        1        ��         ����c   ������������         ����  = >          � g              �  �	        1       ��         ����c   ������������         ����  ? @          � j              �  �	        1       ��         ����c   ������������         ����  A B          � m              
  
        1       ��        ����c   ������������         ����  C D          � p              (  P
        1       ��        ����c   ������������         ����  E F          � s              F  �
        1       ��        ����c   ������������         ����  G H          � v              d  �
        1       ��        ����c   ������������         ����  I J          � y              �          1       ��        ����c   ������������         ����  K L          � |              �  @        1       ��        ����c   ������������         ����  M N          �               �  |        1	       ��        ����c   ������������         ����  & '          y � Fb         >I  �%   	   <      
  ��!        ����
 � �����  �           ����  ( )          ~ � Mf       /  jJ  �2      <     
  ��!        ����
 � �����  �           ����  * +          � � Tj       P  �K  r?      <     
  ��!        ����
 � �����  �           ����  , -          � � [n       q  �L  VL      <     
  ��!       ����
 � �����  �           ����  . /          � � br       �  �M  :Y      <     
  ��!       ����
 � �����  �           ����  0 1          � � iv       �  O  f      <     
  ��!       ����
 � �����  �           ����  3 4          � � pz       �  FP  s      <     
  ��!       ����
 � �����  �           ����  5 6          � � w~       �  rQ  �   ��  <     
  ��!       ����
 � �����  �           ����  7 8          � � ~�       	  �R  ʌ   ��  <     
  ��!       ����
 � �����  �           ����  9 :          � � ��       7	  �S  ��   ��  <	     
  ��!       ����
 7  �  �           ����  1 2            d �            �  F        B        ��"        ����c   ������������         ����  3 4            g �            �  �	        B       ��"        ����c   ������������         ����  5 6            j �            �  �	        B       ��"        ����c   ������������         ����  7 8            m �            
  
        B       ��"       ����c   ������������         ����  9 :            p �            (  P
        B       ��"       ����c   ������������         ����  ; <            s �            F  �
        B       ��"       ����c   ������������         ����  = >            v �            d  �
        B       ��"       ����c   ������������         ����  ? @            y �            �          B       ��"       ����c   ������������         ����  A B            | �            �  @        B       ��"       ����c   ������������         ����  C D             �            �  |        B	       ��"       ����c   ������������         ����  % &          	[ 	]         >I  �%   	   M      
  ��#        ����
 � �����  �           ����  ' (          _ a       /  jJ  �2      M     
  ��#        ����
 � �����  �           ����  ) *          c e       P  �K  r?      M     
  ��#        ����
 � �����  �           ����  + ,          g i       q  �L  VL      M     
  ��#       ����
 � �����  �           ����  - .          !k !m       �  �M  :Y      M     
  ��#       ����
 � �����  �           ����  / 0          'o 'q       �  O  f      M     
  ��#       ����
 � �����  �           ����  2 3          -s -u       �  FP  s      M     
  ��#       ����
 � �����  �           ����  4 5          3w 3y       �  rQ  �   ��  M     
  ��#       ����
 � �����  �           ����  6 7          9{ 9}       	  �R  ʌ   ��  M     
  ��#       ����
 � �����  �           ����  8 9          ? ?�       7	  �S  ��   ��  M	     
  ��#       ����
 7  �  �           ����  0 1          �   �            �  F        S        ��$        ����c   ������������         ����  2 3          �   �            �  �	        S       ��$        ����c   ������������         ����  4 5          �   �            �  �	        S       ��$        ����c   ������������         ����  6 7          �   �            
  
        S       ��$       ����c   ������������         ����  8 9          �   �            (  P
        S       ��$       ����c   ������������         ����  : ;          �   �            F  �
        S       ��$       ����c   ������������         ����  < =          �   �            d  �
        S       ��$       ����c   ������������         ����  > ?          �   �            �          S       ��$       ����c   ������������         ����  @ A          �   �            �  @        S       ��$       ����c   ������������         ����  B C          �   �            �  |        S	       ��$       ����c   ������������         ����� ��                           �����  �s        c      ��9 ��%        ����c �����������������        ����              3 b � /       �  �  ֵ       W        ��&        ���� � ������������         ����              7 f � 2       �  �  º       W       ��&        ���� � ������������         ����              ; j � 5       �  b  ��       W       ��&        ���� � ������������         ����              ? n � 8       �    ��       W       ��&       ���� � ������������         ����              C r � ;         �  ��       W       ��&       ���� � ������������         ����              G v � >         ~  r�       W       ��&       ���� � ������������         ����              K z � A         2  ^�       W       ��&       ���� � ������������         ����               O ~ � D       )  �  J�    	   W       ��&       ���� � ������������         ����   ! "          S � � G       6  �  6�       W       ��&       ���� � ������������         ����   # $          W � � J       B  N   "�       W	       ��&       ���� � ������������         ����              C q � 5       �  #  �      X        ��'        ���� � �����  �           ����              G v � 9       �  �#  �      X       ��'        ���� � �����  �           ����              K { � =       �  �$  &      X       ��'        ���� � �����  �           ����              O � � A         �%  �,      X       ��'       ���� � �����  �           ����              S � � E         f&  03      X       ��'       ���� � �����  �           ����              W � I       #  8'  �9   	   X       ��'       ���� � �����  �           ����     !          [ � M       4  
(  P@      X       ��'       ���� � �����  �           ����   " #          _ � Q       D  �(  �F      X       ��'       ���� � �����  �           ����   $ %          c � U       U  �)  pM      X       ��'       ���� � �����  �           ����   & '          g � Y       f  �*   T      X	       ��'       ���� � �����  �           ����              S � E         �-  �      Y        ��(        ���� � �����  �           ����              W � I       4  �.  x�      Y       ��(        ���� � �����  �           ����              [ � M       J  �/  �      Y       ��(        ���� � �����  �           ����              _ � Q       _  �0  X�   	   Y       ��(       ���� � �����  �           ����               c �  U       u  �1  Ƚ      Y       ��(       ���� � �����  �           ����   ! "          g � 'Y       �  x2  8�      Y       ��(       ���� � �����  �           ����   # $          k � .]       �  h3  ��      Y       ��(       ���� � �����  �           ����   % &          o � 5a       �  X4  �      Y       ��(       ���� � �����  �           ����   ' (          s � <e       �  H5  ��      Y       ��(       ���� � �����  �           ����   ) *          w � Ci       �  86  ��      Y	       ��(       ���� � -  �  �           ����              b � -T       �  �9  �C      Z      	  ��)        ����	 � �����  �           ����              f � 4X       �  ;  <N   
   Z     	  ��)        ����	 � �����  �           ����              j � ;\         <  �X      Z     	  ��)        ����	 � �����  �           ����     !          n � B`         "=  Tc      Z     	  ��)       ����	 � �����  �           ����   " #          r � Id       8  0>  �m      Z     	  ��)       ����	 � �����  �           ����   $ %          v � Ph       S  >?  lx      Z     	  ��)       ����	 � �����  �           ����   & '          z � Wl       n  L@  ��      Z     	  ��)       ����	 � �����  �           ����   ( )          ~ � ^p       �  ZA  ��      Z     	  ��)       ����	 � �����  �           ����   * +          � � et       �  hB  �       Z     	  ��)       ����	 � �����  �           ����   , -          � � lx       �  vC  ��   ��  Z	     	  ��)       ����	 � 7  �  �           ����              q � Uc       �  �G  z   	   [      
  ��*        ����
 � �����  �           ����               v � \g         �H  ^!      [     
  ��*        ����
 � �����  �           ����   ! "          { � ck       $  J  B.      [     
  ��*        ����
 � �����  �           ����   # $          � � jo       E  2K  &;      [     
  ��*       ����
 � �����  �           ����   % &          � � qs       f  ^L  
H      [     
  ��*       ����
 � �����  �           ����   ' (          � � xw       �  �M  �T      [     
  ��*       ����
 � �����  �           ����   ) *          � � {       �  �N  �a      [     
  ��*       ����
 � �����  �           ����   + ,          � � �       �  �O  �n   ��  [     
  ��*       ����
 � �����  �           ����   - .          � � ��       �  Q  �{   ��  [     
  ��*       ����
 � �����  �           ����   / 0          � � ��       	  :R  ~�   ��  [	     
  ��*       ����
 7  �  �            ����             * Y � &       �    *�       �        ��+        ���� � ������������         ����             . ] � )       �  �  �       �       ��+        ���� � ������������         ����             2 a � ,       �  n  �       �       ��+        ���� � ������������         ����             6 e � /       �  "  �       �       ��+       ���� � ������������         ����             : i � 2       �  �  ڻ       �       ��+       ���� � ������������         ����             > m � 5       �  �  ��       �       ��+       ���� � ������������         ����             B q � 8       �  >  ��       �       ��+       ���� � ������������         ����             F u � ;         �  ��    	   �       ��+       ���� � ������������         ����    !          J y � >         �  ��       �       ��+       ���� � ������������         ����  " #          N } � A         Z  v�       �	       ��+       ���� � ������������         ����             : h � ,       �  *!  P	      �        ��,        ���� � �����  �           ����             > m � 0       �  �!  �      �       ��,        ���� � �����  �           ����             B r � 4       �  �"  p      �       ��,        ���� � �����  �           ����             F w � 8       �  �#         �       ��,       ���� � �����  �           ����             J | � <       �  r$  �#      �       ��,       ���� � �����  �           ����             N � � @       �  D%   *   	   �       ��,       ���� � �����  �           ����              R � � D         &  �0      �       ��,       ���� � �����  �           ����  ! "          V � H         �&  @7      �       ��,       ���� � �����  �           ����  # $          Z � L       -  �'  �=      �       ��,       ���� � �����  �           ����  % &          ^ � P       >  �(  `D      �	       ��,       ���� � �����  �           ����             J � � <       �  �+  t�      �        ��-        ���� � �����  �           ����             N � @         �,  �      �       ��-        ���� � �����  �           ����             R � 	D         �-  T�      �       ��-        ���� � �����  �           ����             V � H       2  �.  ģ   	   �       ��-       ���� � �����  �           ����             Z � L       H  �/  4�      �       ��-       ���� � �����  �           ����    !          ^ � P       ]  �0  ��      �       ��-       ���� � �����  �           ����  " #          b � %T       s  t1  �      �       ��-       ���� � �����  �           ����  $ %          f � ,X       �  d2  ��      �       ��-       ���� � �����  �           ����  & '          j � 3\       �  T3  ��      �       ��-       ���� � �����  �           ����  ( )          n � :`       �  D4  d�      �	       ��-       ���� � -  �  �           ����             Y � $K       �  8  (0      �      	  ��.        ����	 � �����  �           ����             ] � +O       �  9  �:   
   �     	  ��.        ����	 � �����  �           ����             a � 2S       �   :  @E      �     	  ��.        ����	 � �����  �           ����              e � 9W       �  .;  �O      �     	  ��.       ����	 � �����  �           ����  ! "          i � @[         <<  XZ      �     	  ��.       ����	 � �����  �           ����  # $          m � G_       !  J=  �d      �     	  ��.       ����	 � �����  �           ����  % &          q � Nc       <  X>  po      �     	  ��.       ����	 � �����  �           ����  ' (          u � Ug       W  f?  �y      �     	  ��.       ����	 � �����  �           ����  ) *          y � \k       r  t@  ��       �     	  ��.       ����	 � �����  �           ����  + ,          } � co       �  �A  �   ��  �	     	  ��.       ����	 � 7  �  �           ����             h � LZ       �  �E  ��   	   �      
  ��/        ����
 � �����  �           ����             m � S^       �  �F  �      �     
  ��/        ����
 � �����  �           ����    !          r � Zb       �  H  �      �     
  ��/        ����
 � �����  �           ����  " #          w � af         >I  �%      �     
  ��/       ����
 � �����  �           ����  $ %          | � hj       /  jJ  �2      �     
  ��/       ����
 � �����  �           ����  & '          � � on       P  �K  r?      �     
  ��/       ����
 � �����  �           ����  ( )          � � vr       q  �L  VL      �     
  ��/       ����
 � �����  �           ����  * +          � � }v       �  �M  :Y   ��  �     
  ��/       ����
 � �����  �           ����  , -          � � �z       �  O  f   ��  �     
  ��/       ����
 � �����  �           ����  . /          � � �~       �  FP  s   ��  �	     
  ��/       ����
 7  �  �           ����             < d � /       �  �  n�       (        ��0        ���� � ������������         ����             @ h � 2       �  V  Z�       (       ��0        ���� � ������������         ����             D l � 5       �  
  F�       (       ��0        ���� � ������������         ����             H p � 8       �  �  2�       (       ��0       ���� � ������������         ����             L t � ;       �  r  �       (       ��0       ���� � ������������         ����             P x � >       �  &  
�       (       ��0       ���� � ������������         ����             T | � A       �  �  ��       (       ��0       ���� � ������������         ����             X � � D       �  �  ��    	   (       ��0       ���� � ������������         ����    !          \ � � G         B  ��       (       ��0       ���� � ������������         ����  " #          ` � � J         �  ��       (	       ��0       ���� � ������������         ����             L s � 5       �  �   0      )        ��1        ���� � �����  �           ����             P x � 9       �  �!  �      )       ��1        ���� � �����  �           ����             T } � =       �  j"  P      )       ��1        ���� � �����  �           ����             X � � A       �  <#  �      )       ��1       ���� � �����  �           ����             \ � � E       �  $  p       )       ��1       ���� � �����  �           ����             ` � � I       �  �$   '   	   )       ��1       ���� � �����  �           ����              d � M         �%  �-      )       ��1       ���� � �����  �           ����  ! "          h � Q         �&   4      )       ��1       ���� � �����  �           ����  # $          l � U       %  V'  �:      )       ��1       ���� � �����  �           ����  % &          p � Y       6  ((  @A      )	       ��1       ���� � �����  �           ����             \ � � E       �  p+  ��      *        ��2        ���� � �����  �           ����             ` � I       �  `,  `�      *       ��2        ���� � �����  �           ����             d � M         P-  З      *       ��2        ���� � �����  �           ����             h � Q       )  @.  @�   	   *       ��2       ���� � �����  �           ����             l � U       ?  0/  ��      *       ��2       ���� � �����  �           ����    !          p � !Y       T   0   �      *       ��2       ���� � �����  �           ����  " #          t � (]       j  1  ��      *       ��2       ���� � �����  �           ����  $ %          x � /a       �   2   �      *       ��2       ���� � �����  �           ����  & '          | � 6e       �  �2  p�      *       ��2       ���� � �����  �           ����  ( )          � � =i       �  �3  ��      *	       ��2       ���� � -  �  �           ����             k � 'T       �  �7  @,      +      	  ��3        ����	 � �����  �           ����             o � .X       �  �8  �6   
   +     	  ��3        ����	 � �����  �           ����             s � 5\       �  �9  XA      +     	  ��3        ����	 � �����  �           ����              w � <`       �  �:  �K      +     	  ��3       ����	 � �����  �           ����  ! "          { � Cd       �  �;  pV      +     	  ��3       ����	 � �����  �           ����  # $           � Jh         �<  �`      +     	  ��3       ����	 � �����  �           ����  % &          � � Ql       2  �=  �k      +     	  ��3       ����	 � �����  �           ����  ' (          � � Xp       M  ?  v      +     	  ��3       ����	 � �����  �           ����  ) *          � � _t       h  @  ��       +     	  ��3       ����	 � �����  �           ����  + ,          � � fx       �  A  ,�   ��  +	     	  ��3       ����	 � 7  �  �           ����             z � Oc       �  VE  ��   	   ,      
  ��4        ����
 � �����  �           ����              � Vg       �  �F  �      ,     
  ��4        ����
 � �����  �           ����    !          � � ]k       �  �G  z      ,     
  ��4        ����
 � �����  �           ����  " #          � � do         �H  ^!      ,     
  ��4       ����
 � �����  �           ����  $ %          � � ks       $  J  B.      ,     
  ��4       ����
 � �����  �           ����  & '          � � rw       E  2K  &;      ,     
  ��4       ����
 � �����  �           ����  ( )          � � y{       f  ^L  
H      ,     
  ��4       ����
 � �����  �           ����  * +          � � �       �  �M  �T   ��  ,     
  ��4       ����
 � �����  �           ����  , -          � � ��       �  �N  �a   ��  ,     
  ��4       ����
 � �����  �           ����  . /          � � ��       �  �O  �n   ��  ,	     
  ��4       ����
 7  �  �            ����             ' V � #       %  �  ��       �        ��5        ���� � ������������         ����             + Z � &       2  ^  ��       �       ��5        ���� � ������������         ����             / ^ � )       >     ~�       �       ��5        ���� � ������������         ����             3 b � ,       K  �   j�       �       ��5       ���� � ������������         ����             7 f � /       W  z!  V�       �       ��5       ���� � ������������         ����             ; j � 2       d  ."  B�       �       ��5       ���� � ������������         ����             ? n � 5       q  �"  .�       �       ��5       ���� � ������������         ����             C r � 8       }  �#  �    	   �       ��5       ���� � ������������         ����    !          G v � ;       �  J$  �       �       ��5       ���� � ������������         ����  " #          K z � >       �  �$  �      �	       ��5       ���� � ������������         ����             7 e � )       /  �'  p>      �        ��6        ���� � �����  �            ����             ; j � -       @  �(   E      �       ��6        ���� � �����  �            ����             ? o � 1       P  r)  �K      �       ��6        ���� � �����  �            ����             C t � 5       a  D*   R      �       ��6       ���� � �����  �            ����             G y � 9       r  +  �X      �       ��6       ���� � �����  �            ����             K ~ � =       �  �+  @_   	   �       ��6       ���� � �����  �            ����              O � � A       �  �,  �e      �       ��6       ���� � �����  �            ����  ! "          S � E       �  �-  `l      �       ��6       ���� � �����  �            ����  # $          W � I       �  ^.  �r      �       ��6       ���� � �����  �            ����  % &          [ � M       �  0/  �y      �	       ��6       ���� � �����  �            ����             G } � 9       �  x2  8�      �        ��7        ���� � �����  �  !         ����             K � � =       �  h3  ��      �       ��7        ���� � �����  �  !         ����             O � A       �  X4  �      �       ��7        ���� � �����  �  !         ����             S � E       �  H5  ��   	   �       ��7       ���� � �����  �  !         ����             W � I       �  86  ��      �       ��7       ���� � �����  �  !         ����    !          [ � M       �  (7  h�      �       ��7       ���� � �����  �  !         ����  " #          _ � "Q         8  ��      �       ��7       ���� � �����  �  !         ����  $ %          c � )U       "  9  H      �       ��7       ���� � �����  �  !         ����  & '          g � 0Y       7  �9  �	      �       ��7       ���� � �����  �  !         ����  ( )          k � 7]       M  �:  (      �	       ��7       ���� � -  �  �  !         ����             V � !H       D  �>  �r      �      	  ��8        ����	 � �����  �  "         ����             Z � (L       _  �?  }   
   �     	  ��8        ����	 � �����  �  "         ����             ^ � /P       z  �@  ��      �     	  ��8        ����	 � �����  �  "         ����              b � 6T       �  �A  4�      �     	  ��8       ����	 � �����  �  "         ����  ! "          f � =X       �  �B  ��      �     	  ��8       ����	 � �����  �  "         ����  # $          j � D\       �  �C  L�      �     	  ��8       ����	 � �����  �  "         ����  % &          n � K`       �  �D  ر      �     	  ��8       ����	 � �����  �  "         ����  ' (          r � Rd         
F  d�      �     	  ��8       ����	 � �����  �  "         ����  ) *          v � Yh         G  ��       �     	  ��8       ����	 � �����  �  "         ����  + ,          z � `l       7  &H  |�   ��  �	     	  ��8       ����	 � 7  �  �  "         ����             e � IW       f  ^L  
H   	   �      
  ��9        ����
 � �����  �  #         ����             j � P[       �  �M  �T      �     
  ��9        ����
 � �����  �  #         ����    !          o � W_       �  �N  �a      �     
  ��9        ����
 � �����  �  #         ����  " #          t � ^c       �  �O  �n      �     
  ��9       ����
 � �����  �  #         ����  $ %          y � eg       �  Q  �{      �     
  ��9       ����
 � �����  �  #         ����  & '          ~ � lk       	  :R  ~�      �     
  ��9       ����
 � �����  �  #         ����  ( )          � � so       ,	  fS  b�      �     
  ��9       ����
 � �����  �  #         ����  * +          � � zs       M	  �T  F�   ��  �     
  ��9       ����
 � �����  �  #         ����  , -          � � �w       n	  �U  *�   ��  �     
  ��9       ����
 � �����  �  #         ����  . /          � � �{       �	  �V  �   ��  �	     
  ��9       ����
 7  �  �  #         ����             B q � >       	    ��       �        ��:        ���� � ������������$         ����             F u � A         �  ��       �       ��:        ���� � ������������$         ����             J y � D       "  �  ��       �       ��:        ���� � ������������$         ����             N } � G       /  6  z�       �       ��:       ���� � ������������$         ����             R � � J       ;  �  f�       �       ��:       ���� � ������������$         ����             V � � M       H  �   R�       �       ��:       ���� � ������������$         ����             Z � � P       U  R!  >�       �       ��:       ���� � ������������$         ����              ^ � � S       a  "  *�    	   �       ��:       ���� � ������������$         ����  ! "          b � V       n  �"  �       �       ��:       ���� � ������������$         ����  # $          f � Y       z  n#  �       �	       ��:       ���� � ������������$         ����             R � � D         >&  �1      �        ��;        ���� � �����  �  %         ����             V � � H          '  �8      �       ��;        ���� � �����  �  %         ����             Z � � L       0  �'  ?      �       ��;        ���� � �����  �  %         ����             ^ � P       A  �(  �E      �       ��;       ���� � �����  �  %         ����             b � T       R  �)  0L      �       ��;       ���� � �����  �  %         ����             f � X       c  X*  �R   	   �       ��;       ���� � �����  �  %         ����    !          j � \       t  *+  PY      �       ��;       ���� � �����  �  %         ����  " #          n � `       �  �+  �_      �       ��;       ���� � �����  �  %         ����  $ %          r � #d       �  �,  pf      �       ��;       ���� � �����  �  %         ����  & '          v � )h       �  �-   m      �	       ��;       ���� � �����  �  %         ����             b � T       f  �0  (�      �        ��<        ���� � �����  �  &         ����             f � X       |  �1  ��      �       ��<        ���� � �����  �  &         ����             j � !\       �  �2  �      �       ��<        ���� � �����  �  &         ����             n � (`       �  �3  x�   	   �       ��<       ���� � �����  �  &         ����              r � /d       �  �4  ��      �       ��<       ���� � �����  �  &         ����  ! "          v � 6h       �  �5  X�      �       ��<       ���� � �����  �  &         ����  # $          z � =l       �  �6  ��      �       ��<       ���� � �����  �  &         ����  % &          ~ � Dp       �  x7  8�      �       ��<       ���� � �����  �  &         ����  ' (          � � Kt         h8  ��      �       ��<       ���� � �����  �  &         ����  ) *          � � Rx       )  X9        �	       ��<       ���� � -  �  �  &         ����             q � <c         =  �b      �        ��=        ����	 � �����  �  '         ����             u � Cg       7  &>  |m   
   �       ��=        ����	 � �����  �  '         ����             y � Jk       R  4?  x      �       ��=        ����	 � �����  �  '         ����    !          } � Qo       m  B@  ��      �       ��=       ����	 � �����  �  '         ����  " #          � � Xs       �  PA   �      �       ��=       ����	 � �����  �  '         ����  $ %          � � _w       �  ^B  ��      �       ��=       ����	 � �����  �  '         ����  & '          � � f{       �  lC  8�      �       ��=       ����	 � �����  �  '         ����  ( )          � � m       �  zD  Ĭ      �       ��=       ����	 � �����  �  '         ����  * +          � � t�       �  �E  P�       �       ��=       ����	 � �����  �  '         ����  , -          � � {�         �F  ��   ��  �	       ��=       ����	 � 7  �  �  '         ����             � � dr       :  �J  �6   	   �      	  ��>        ����
 � �����  �  (         ����              � � kv       [  �K  �C      �     	  ��>        ����
 � �����  �  (         ����  ! "          � � rz       |  &M  �P      �     	  ��>        ����
 � �����  �  (         ����  # $          � � y~       �  RN  �]      �     	  ��>       ����
 � �����  �  (         ����  % &          � � ��       �  ~O  jj      �     	  ��>       ����
 � �����  �  (         ����  ' (          � � ��       �  �P  Nw      �     	  ��>       ����
 � �����  �  (         ����  ) *          � � ��        	  �Q  2�      �     	  ��>       ����
 � �����  �  (         ����  + ,          � � ��       !	  S  �   ��  �     	  ��>       ����
 � �����  �  (         ����  - .          � � ��       B	  .T  ��   ��  �     	  ��>       ����
 � �����  �  (         ����  / 0          � � ��       c	  ZU  ު   ��  �	     	  ��>       ����
 7  �  �  (          ����             9 h � 5       �  �  ��       Z        ��?        ���� � ������������)         ����             = l � 8       �  >  ��       Z       ��?        ���� � ������������)         ����             A p � ;         �  ��       Z       ��?        ���� � ������������)         ����             E t � >         �  ��       Z       ��?       ���� � ������������)         ����             I x � A         Z  v�       Z       ��?       ���� � ������������)         ����             M | � D       ,    b�       Z       ��?       ���� � ������������)         ����             Q � � G       9  �  N�       Z       ��?       ���� � ������������)         ����             U � � J       E  v   :�    	   Z       ��?       ���� � ������������)         ����    !          Y � � M       R  *!  &�       Z       ��?       ���� � ������������)         ����  " #          ] � � P       ^  �!  �       Z	       ��?       ���� � ������������)         ����             I w � ;       �  �$  p%      [        ��@        ���� � �����  �  *         ����             M | � ?          �%   ,      [       ��@        ���� � �����  �  *         ����             Q � � C         R&  �2      [       ��@        ���� � �����  �  *         ����             U � � G       !  $'   9      [       ��@       ���� � �����  �  *         ����             Y � K       2  �'  �?      [       ��@       ���� � �����  �  *         ����             ] � O       C  �(  @F   	   [       ��@       ���� � �����  �  *         ����              a � S       T  �)  �L      [       ��@       ���� � �����  �  *         ����  ! "          e � W       d  l*  `S      [       ��@       ���� � �����  �  *         ����  # $          i � [       u  >+  �Y      [       ��@       ���� � �����  �  *         ����  % &          m �  _       �  ,  �`      [	       ��@       ���� � �����  �  *         ����             Y � 
K       B  X/  �      \        ��A        ���� � �����  �  +         ����             ] � O       X  H0  ��      \       ��A        ���� � �����  �  +         ����             a � S       n  81  ��      \       ��A        ���� � �����  �  +         ����             e � W       �  (2  h�   	   \       ��A       ���� � �����  �  +         ����             i � &[       �  3  ��      \       ��A       ���� � �����  �  +         ����    !          m � -_       �  4  H�      \       ��A       ���� � �����  �  +         ����  " #          q � 4c       �  �4  ��      \       ��A       ���� � �����  �  +         ����  $ %          u � ;g       �  �5  (�      \       ��A       ���� � �����  �  +         ����  & '          y � Bk       �  �6  ��      \       ��A       ���� � �����  �  +         ����  ( )          } � Io         �7  �      \	       ��A       ���� � -  �  �  +         ����             h � 3Z       �  �;  PS      ]      	  ��B        ����	 � �����  �  ,         ����             l � :^         �<  �]   
   ]     	  ��B        ����	 � �����  �  ,         ����             p � Ab       *  �=  hh      ]     	  ��B        ����	 � �����  �  ,         ����              t � Hf       E  �>  �r      ]     	  ��B       ����	 � �����  �  ,         ����  ! "          x � Oj       `  �?  �}      ]     	  ��B       ����	 � �����  �  ,         ����  # $          | � Vn       {  �@  �      ]     	  ��B       ����	 � �����  �  ,         ����  % &          � � ]r       �  �A  ��      ]     	  ��B       ����	 � �����  �  ,         ����  ' (          � � dv       �  �B  $�      ]     	  ��B       ����	 � �����  �  ,         ����  ) *          � � kz       �  �C  ��       ]     	  ��B       ����	 � �����  �  ,         ����  + ,          � � r~       �  E  <�   ��  ]	     	  ��B       ����	 � 7  �  �  ,         ����             w � [i         >I  �%   	   ^      
  ��C        ����
 � �����  �  -         ����             | � bm       /  jJ  �2      ^     
  ��C        ����
 � �����  �  -         ����    !          � � iq       P  �K  r?      ^     
  ��C        ����
 � �����  �  -         ����  " #          � � pu       q  �L  VL      ^     
  ��C       ����
 � �����  �  -         ����  $ %          � � wy       �  �M  :Y      ^     
  ��C       ����
 � �����  �  -         ����  & '          � � ~}       �  O  f      ^     
  ��C       ����
 � �����  �  -         ����  ( )          � � ��       �  FP  s      ^     
  ��C       ����
 � �����  �  -         ����  * +          � � ��       �  rQ  �   ��  ^     
  ��C       ����
 � �����  �  -         ����  , -          � � ��       	  �R  ʌ   ��  ^     
  ��C       ����
 � �����  �  -         ����  . /          � � ��       7	  �S  ��   ��  ^	     
  ��C       ����
 7  �  �  -            ��              ( + 4 .      �����
  �         �       �    D        ���� � ������������.            ��              * . 9 0      ����          �      �    D        ���� � ������������.            ��              , 1 > 2      ����,  X        �      �    D        ���� � ������������.            ��   	           . 4 C 4      ����J  �        �      �    D        ���� � ������������.            ��  
            0 7 H 6      ����h  �        �      �    D        ���� � ������������.            ��              2 : M 8      �����          �      �    D        ���� � ������������.            ��              4 = R :      �����  H        �      �    D        ���� � ������������.            ��              6 @ W <      �����  �        �      �    D        ���� � ������������.            ��              8 C \ >      �����  �        �      �    D        ���� � ������������.            ��              : F a @      �����  �        � 	     �    D        ���� � ������������.           ��              * 3 O 0 (     ����v  b%        �       �    E        ���� � ������������/           ��              - 6 T 2 (     �����  &        �      �    E        ���� � ������������/           ��  	 
           0 9 Y 4 (     �����  �&        �      �    E        ���� � ������������/           ��              3 < ^ 6 (     ����*  ~'        �      �    E        ���� � ������������/           ��              6 ? c 8 (     ����f  2(        �      �    E        ���� � ������������/           ��              9 B h : (     �����  �(        �      �    E        ���� � ������������/           ��              < E m < (     �����  �)        �      �    E        ���� � ������������/           ��              ? H r > (     ����  N*        �      �    E        ���� � ������������/           ��              B K w @ (     ����V  +        �      �    E        ���� � ������������/           ��              E N | B (     �����  �+        � 	     �    E        ���� � ������������/          ��   	           - : i 2 2     �����  >        �       �    F        ���� � ������������0          ��  
            0 > n 5 2     �����  p?        �      �    F        ���� � ������������0          ��              3 B s 8 2     ����6  �@        �      �    F        ���� � ������������0          ��              6 F x ; 2     �����  @B        �      �    F        ���� � ������������0          ��              9 J } > 2     �����  �C        �      �    F        ���� � ������������0          ��              < N � A 2     ����D  E        �      �    F        ���� � ������������0          ��              ? R � D 2     �����  xF        �      �    F        ���� � ������������0          ��              B V � G 2     �����  �G        �      �    F        ���� � ������������0          ��              E Z � J 2     ����R  HI        �      �    F        ���� � ������������0          ��              H ^ � M 2     �����  �J        � 	     �    F        ���� � ������������0         	 ��              5 K � 4 <     ����  dd        �       �    G        ���� � ������������1         	 ��              8 O � 7 <     �����  �f        �      �    G        ���� � ������������1         	 ��              ; S � : <     ����  i        �      �    G        ���� � ������������1         	 ��              > W � = <     ����|  lk        �      �    G        ���� � ������������1         	 ��              A [ � @ <     �����  �m        �      �    G        ���� � ������������1         	 ��              D _ � C <     ����l  p        �      �    G        ���� � ������������1         	 ��              G c � F <     �����  tr        �      �    G        ���� � ������������1         	 ��              J g � I <     ����\  �t        �      �    G        ���� � ������������1         	 ��              M k � L <     �����  $w        �      �    G        ���� � ������������1         	 ��              P o � O <     ����L  |y        � 	     �    G        ���� � ������������1         
 ��              < [ � ; F     ����,  �        �       �    H        ���� � ������������2         
 ��              ? _ � > F     �����  ��        �      �    H        ���� � ������������2         
 ��              B c � A F     ����X  �        �      �    H        ���� � ������������2          ��              E g � D F     �����  ��        �      �    H        ���� � ������������2          ��              H k � G F     �����  �        �      �    H        ���� � ������������2          ��              K o � J F     ����  ��        �      �    H        ���� � ������������2          ��              N s � M F     �����   �        �      �    H        ���� � ������������2          ��              Q w � P F     ����F  ��        �      �    H        ���� � ������������2          ��              T { � S F     �����  (�        �      �    H        ���� � ������������2          ��    !           W  � V F     ����r  ��        � 	     �    H        ���� � ������������2          ��              C j � B P     �����!  ��        �       �    I        ���� � ������������3          ��              G n � E P     ����~"  r�        �      �    I        ���� � ������������3          ��              K r � H P     ����2#  ^�        �      �    I        ���� � ������������3          ��              O v � K P     �����#  J�        �      �    I        ���� � ������������3          ��              S z � N P     �����$  6        �      �    I        ���� � ������������3          ��              W ~ � Q P     ����N%  "       �      �    I        ���� � ������������3          ��              [ � � T P     ����&  
       �      �    I        ���� � ������������3          ��               _ � � W P     �����&  �       �      �    I        ���� � ������������3          ��  ! "           c � � Z P     ����j'  �       �      �    I        ���� � ������������3          ��  # $           g � � ] P     ����(  �       � 	     �    I        ���� � ������������3          ��              S y � H Z     �����*  pW       �       �    J        ���� � �����  �  4          ��              W ~ � L Z     �����+   ^       �      �    J        ���� � �����  �  4          ��              [ � � P Z     �����,  �d       �      �    J        ���� � �����  �  4          ��              _ � � T Z     ����d-   k       �      �    J        ���� � �����  �  4          ��              c � � X Z     ����6.  �q       �      �    J        ���� � �����  �  4          ��              g � \ Z     ����/  @x       �      �    J        ���� � �����  �  4          ��    !           k � ` Z     �����/  �~       �      �    J        ���� � �����  �  4          ��  " #           o � d Z     �����0  `�       �      �    J        ���� � �����  �  4          ��  $ %           s � h Z     ����~1  ��       �      �    J        ���� � �����  �  4          ��  & '           w � l Z     ����P2  ��       � 	     �    J        ���� � �����  �  4          ��              c � X d     �����5  X�       �       �    K        ���� � �����  �  5          ��              g � \ d     �����6  ��       �      �    K        ���� � �����  �  5          ��              k � ` d     ����x7  8�       �      �    K        ���� � �����  �  5          ��              o � d d     ����h8  ��       �      �    K        ���� � �����  �  5          ��               s � #h d     ����X9         �      �    K        ���� � �����  �  5          ��  ! "           w � *l d     ����H:  �       �      �    K        ���� � �����  �  5          ��  # $           { � 1p d     ����8;  �       �      �    K        ���� � �����  �  5          ��  % &            � 8t d     ����(<  h       �      �    K        ���� � �����  �  5          ��  ' (           � � ?x d     ����=  �%       �      �    K        ���� � �����  �  5          ��  ) *           � � F| d     ����>  H.       � 	     �    K        ���� � �����  �  5          ��              r � 0g n     �����A  Б       �       �    L        ����	 � �����  �  6          ��              v � 7k n     �����B  \�       �      �    L        ����	 � �����  �  6          ��              z � >o n     �����C  �       �      �    L        ����	 � �����  �  6          ��    !           ~ � Es n     �����D  t�       �      �    L        ����	 � �����  �  6          ��  " #           � � Lw n     ���� F   �       �      �    L        ����	 � �����  �  6          ��  $ %           � � S{ n     ����G  ��       �      �    L        ����	 � �����  �  6          ��  & '           � � Z n     ����H  �       �      �    L        ����	 � �����  �  6          ��  ( )           � � a� n     ����*I  ��       �      �    L        ����	 � �����  �  6          ��  * +           � � h� n     ����8J  0�       �      �    L        ����	 � �����  �  6          ��  , -           � � o� n     ����FK  ��       � 	     �    L        ����	 � �����  �  6          ����	                        ����  .J       
      �� ��M        ���� � ������������7          ����	                !        ����.  \       
     �� ��M        ���� � ������������7          ����	                &        ����L  �       
     �� ��M        ���� � ������������7          ����	   	             +        ����j  �       
     �� ��M       ���� � ������������7          ����	  
              0        �����         
     �� ��M       ���� � ������������7          ����	               " 5         �����  L       
     �� ��M       ���� � ������������7          ����	               % : "       �����  �       
     �� ��M       ���� � ������������7          ����	               ( ? $       �����  �       
     �� ��M       ���� � ������������7          ����	                + D &       ����           
     �� ��M       ���� � ������������7          ����	              " . I (       ����  <       
	     �� ��M       ���� � ������������7          ����	                7        �����  �.             �� ��N        ���� � ������������8          ����	                <        �����  v/            �� ��N        ���� � ������������8          ����	  	 
            ! A        ����  *0            �� ��N        ���� � ������������8          ����	               $ F        ����J  �0            �� ��N       ���� � ������������8          ����	              ! ' K         �����  �1            �� ��N       ���� � ������������8          ����	              $ * P "       �����  F2            �� ��N       ���� � ������������8          ����	              ' - U $       �����  �2            �� ��N       ���� � ������������8          ����	              * 0 Z &       ����:  �3            �� ��N       ���� � ������������8          ����	              - 3 _ (       ����v  b4            �� ��N       ���� � ������������8          ����	              0 6 d *       �����  5       	     �� ��N       ���� � ������������8         ����	   	            " Q        �����  �J             �� ��O        ���� � ������������9         ����	  
              & V        �����  �K            �� ��O        ���� � ������������9         ����	              # * [         ����V  XM            �� ��O        ���� � ������������9         ����	              & . ` #       �����  �N            �� ��O       ���� � ������������9         ����	              ) 2 e &       ����
  (P            �� ��O       ���� � ������������9         ����	              , 6 j )       ����d  �Q            �� ��O       ���� � ������������9         ����	              / : o ,       �����  �R            �� ��O       ���� � ������������9         ����	              2 > t /       ����  `T            �� ��O       ���� � ������������9         ����	              5 B y 2       ����r  �U            �� ��O       ���� � ������������9         ����	              8 F ~ 5       �����  0W       	     �� ��O       ���� � ������������9         ����	              % 3 j        ����4  t             �� ��P        ���� � ������������:         ����	              ( 7 p !       �����  \v            �� ��P        ���� � ������������:         ����	              + ; v $       ����$  �x            �� ��P        ���� � ������������:         ����	              . ? | '       �����  {            �� ��P       ���� � ������������:         ����	              1 C � *       ����  d}            �� ��P       ���� � ������������:         ����	              4 G � -       �����  �            �� ��P       ���� � ������������:         ����	              7 K � 0       ����  �            �� ��P       ���� � ������������:         ����	              : O � 3       ����|  l�            �� ��P       ���� � ������������:         ����	              = S � 6       �����  Ć            �� ��P       ���� � ������������:         ����	              @ W � 9       ����l  �       	     �� ��P       ���� � ������������:         ����	              , C � %       ����L  ȯ             �� ��Q        ���� � ������������;         ����	              / G � (       �����  L�            �� ��Q        ���� � ������������;         ����	              2 K � +       ����x  ж            �� ��Q        ���� � ������������;         ����	              5 O � .       ����  T�            �� ��Q       ���� � ������������;         ����	              8 S � 1       �����  ؽ            �� ��Q       ���� � ������������;         ����	              ; W � 4       ����:   \�            �� ��Q       ���� � ������������;         ����	              > [ � 7       �����   ��            �� ��Q       ���� � ������������;         ����	              A _ � :       ����f!  d�            �� ��Q       ���� � ������������;         ����	              D c � =       �����!  ��    
        �� ��Q       ���� � ������������;         ����	    !           G g � @       �����"  l�    	   	     �� ��Q       ���� � ������������;         ����	              3 R � ,       �����$  f            �� ��R        ���� � ������������<         ����	              7 V � /       �����%  R           �� ��R        ���� � ������������<         ����	              ; Z � 2       ����R&  >           �� ��R        ���� � ������������<         ����	              ? ^ � 5       ����'  *           �� ��R       ���� � ������������<         ����	              C b � 8       �����'             �� ��R       ���� � ������������<         ����	              G f � ;       ����n(             �� ��R       ���� � ������������<         ����	              K j � >       ����")  �           �� ��R       ���� � ������������<         ����	               O n � A       �����)  �$   	        �� ��R       ���� � ������������<         ����	  ! "           S r � D       �����*  �)           �� ��R       ���� � ������������<         ����	  # $           W v � G       ����>+  �.      	     �� ��R       ���� � ������������<         ����	              C a � 2       ����.  pp            �� ��S        ���� � �����  �  =         ����	              G f � 6       �����.   w           �� ��S        ���� � �����  �  =         ����	              K k � :       �����/  �}           �� ��S        ���� � �����  �  =         ����	              O p � >       �����0   �           �� ��S       ���� � �����  �  =         ����	              S u � B       ����V1  ��           �� ��S       ���� � �����  �  =         ����	              W z � F       ����(2  @�   	        �� ��S       ���� � �����  �  =         ����	    !           [  � J       �����2  З           �� ��S       ���� � �����  �  =         ����	  " #           _ � � N       �����3  `�           �� ��S       ���� � �����  �  =         ����	  $ %           c � � R       �����4  �           �� ��S       ���� � �����  �  =         ����	  & '           g � V       ����p5  ��      	     �� ��S       ���� � �����  �  =         ����	              S y � B       �����8  x�            �� ��T        ���� � �����  �  >         ����	              W ~ � F       �����9  �           �� ��T        ���� � �����  �  >         ����	              [ � � J       �����:  X           �� ��T        ���� � �����  �  >         ����	              _ � N       �����;  �   	        �� ��T       ���� � �����  �  >         ����	               c � R       ����x<  8            �� ��T       ���� � �����  �  >         ����	  ! "           g � V       ����h=  �(           �� ��T       ���� � �����  �  >         ����	  # $           k � Z       ����X>  1           �� ��T       ���� � �����  �  >         ����	  % &           o �  ^       ����H?  �9           �� ��T       ���� � �����  �  >         ����	  ' (           s � 'b       ����8@  �A           �� ��T       ���� � �����  �  >         ����	  ) *           w � .f       ����(A  hJ      	     �� ��T       ���� � �����  �  >         ����	              b � Q       �����D  �            �� ��U        ����	 � �����  �  ?         ����	              f � U       �����E  ��   
        �� ��U        ����	 � �����  �  ?         ����	              j � &Y       ����G  (�           �� ��U        ����	 � �����  �  ?         ����	    !           n � -]       ����H  ��           �� ��U       ����	 � �����  �  ?         ����	  " #           r � 4a       ���� I  @�           �� ��U       ����	 � �����  �  ?         ����	  $ %           v � ;e       ����.J  ��           �� ��U       ����	 � �����  �  ?         ����	  & '           z � Bi       ����<K  X�           �� ��U       ����	 � �����  �  ?         ����	  ( )           ~ � Im       ����JL  ��           �� ��U       ����	 � �����  �  ?         ����	  * +           � � Pq       ����XM  p            �� ��U       ����	 � �����  �  ?         ����	  , -           � � Wu       ����fN  �   ��  	     �� ��U       ����	 � �����  �  ?          ����
                %        �����  t1       d      �� ��V        ���� � ������������@          ����
                * !       �����  <       d     �� ��V        ���� � ������������@          ����
               " / #       �����  x       d     �� ��V        ���� � ������������@          ����
   	            % 4 %       �����  �       d     �� ��V       ���� � ������������@          ����
  
            ! ( 9 '       �����  �       d     �� ��V       ���� � ������������@          ����
              # + > )       ����  ,       d     �� ��V       ���� � ������������@          ����
              % . C +       ����4  h       d     �� ��V       ���� � ������������@          ����
              ' 1 H -       ����R  �       d     �� ��V       ���� � ������������@          ����
              ) 4 M /       ����p  �       d     �� ��V       ���� � ������������@          ����
              + 7 R 1       �����         d	     �� ��V       ���� � ������������@          ����
               $ @ !       ����  *       e      �� ��W        ���� � ������������A          ����
               ' E #       ����B  �*       e     �� ��W        ���� � ������������A          ����
  	 
           " * J %       ����~  z+       e     �� ��W        ���� � ������������A          ����
              % - O '       �����  .,       e     �� ��W       ���� � ������������A          ����
              ( 0 T )       �����  �,       e     �� ��W       ���� � ������������A          ����
              + 3 Y +       ����2  �-       e     �� ��W       ���� � ������������A          ����
              . 6 ^ -       ����n  J.       e     �� ��W       ���� � ������������A          ����
              1 9 c /       �����  �.       e     �� ��W       ���� � ������������A          ����
              4 < h 1       �����  �/       e     �� ��W       ���� � ������������A          ����
              7 ? m 3       ����"  f0       e	     �� ��W       ���� � ������������A         ����
   	           $ + Z #       ����  HD       f      �� ��X        ���� � ������������B         ����
  
            ' / _ &       ����l  �E       f     �� ��X        ���� � ������������B         ����
              * 3 d )       �����  G       f     �� ��X        ���� � ������������B         ����
              - 7 i ,       ����   �H       f     �� ��X       ���� � ������������B         ����
              0 ; n /       ����z  �I       f     �� ��X       ���� � ������������B         ����
              3 ? s 2       �����  PK       f     �� ��X       ���� � ������������B         ����
              6 C x 5       ����.  �L       f     �� ��X       ���� � ������������B         ����
              9 G } 8       �����   N       f     �� ��X       ���� � ������������B         ����
              < K � ;       �����  �O       f     �� ��X       ���� � ������������B         ����
              ? O � >       ����<  �P       f	     �� ��X       ���� � ������������B         ����
              , < s '       �����  4l       g      �� ��Y        ���� � ������������C         ����
              / @ y *       ����  �n       g     �� ��Y        ���� � ������������C         ����
              2 D  -       �����  �p       g     �� ��Y        ���� � ������������C         ����
              5 H � 0       ����  <s       g     �� ��Y       ���� � ������������C         ����
              8 L � 3       �����  �u       g     �� ��Y       ���� � ������������C         ����
              ; P � 6       �����  �w       g     �� ��Y       ���� � ������������C         ����
              > T � 9       ����t  Dz       g     �� ��Y       ���� � ������������C         ����
              A X � <       �����  �|       g     �� ��Y       ���� � ������������C         ����
              D \ � ?       ����d  �~       g     �� ��Y       ���� � ������������C         ����
              G ` � B       �����  L�       g	     �� ��Y       ���� � ������������C         ����
              3 L � .       �����  h�       h      �� ��Z        ���� � ������������D         ����
              6 P � 1       ����R  �       h     �� ��Z        ���� � ������������D         ����
              9 T � 4       �����  p�       h     �� ��Z        ���� � ������������D         ����
              < X � 7       ����~  ��       h     �� ��Z       ���� � ������������D         ����
              ? \ � :       ����  x�       h     �� ��Z       ���� � ������������D         ����
              B ` � =       �����  ��       h     �� ��Z       ���� � ������������D         ����
              E d � @       ����@  ��       h     �� ��Z       ���� � ������������D         ����
              H h � C       �����  �       h     �� ��Z       ���� � ������������D         ����
              K l � F       ����l   ��    
   h     �� ��Z       ���� � ������������D         ����
    !           N p � I       ����!  �    	   h	     �� ��Z       ���� � ������������D         ����
              : [ � 5       ����Z#  v�       i      �� ��[        ���� � ������������E         ����
              > _ � 8       ����$  b�       i     �� ��[        ���� � ������������E         ����
              B c � ;       �����$  N      i     �� ��[        ���� � ������������E         ����
              F g � >       ����v%  :      i     �� ��[       ���� � ������������E         ����
              J k � A       ����*&  &      i     �� ��[       ���� � ������������E         ����
              N o � D       �����&        i     �� ��[       ���� � ������������E         ����
              R s � G       �����'  �      i     �� ��[       ���� � ������������E         ����
               V w � J       ����F(  �   	   i     �� ��[       ���� � ������������E         ����
  ! "           Z { � M       �����(  �      i     �� ��[       ���� � ������������E         ����
  # $           ^  � P       �����)  �#      i	     �� ��[       ���� � ������������E         ����
              J j � ;       ����~,  �c      j      �� ��\        ���� � �����  �  F         ����
              N o � ?       ����P-  �j      j     �� ��\        ���� � �����  �  F         ����
              R t � C       ����".  q      j     �� ��\        ���� � �����  �  F         ����
              V y � G       �����.  �w      j     �� ��\       ���� � �����  �  F         ����
              Z ~ � K       �����/  0~      j     �� ��\       ���� � �����  �  F         ����
              ^ � � O       �����0  ��   	   j     �� ��\       ���� � �����  �  F         ����
    !           b � � S       ����j1  P�      j     �� ��\       ���� � �����  �  F         ����
  " #           f � W       ����<2  ��      j     �� ��\       ���� � �����  �  F         ����
  $ %           j � [       ����3  p�      j     �� ��\       ���� � �����  �  F         ����
  & '           n � _       �����3   �      j	     �� ��\       ���� � �����  �  F         ����
              Z � � K       ����(7  h�      k      �� ��]        ���� � �����  �  G         ����
              ^ � � O       ����8  ��      k     �� ��]        ���� � �����  �  G         ����
              b � S       ����9  H      k     �� ��]        ���� � �����  �  G         ����
              f � W       �����9  �	   	   k     �� ��]       ���� � �����  �  G         ����
               j � [       �����:  (      k     �� ��]       ���� � �����  �  G         ����
  ! "           n � _       �����;  �      k     �� ��]       ���� � �����  �  G         ����
  # $           r � "c       �����<  #      k     �� ��]       ���� � �����  �  G         ����
  % &           v � )g       �����=  x+      k     �� ��]       ���� � �����  �  G         ����
  ' (           z � 0k       �����>  �3      k     �� ��]       ���� � �����  �  G         ����
  ) *           ~ � 7o       �����?  X<      k	     �� ��]       ���� � �����  �  G         ����
              i � !Z       ����XC  p�      l      �� ��^        ����	 � �����  �  H         ����
              m � (^       ����fD  ��   
   l     �� ��^        ����	 � �����  �  H         ����
              q � /b       ����tE  ��      l     �� ��^        ����	 � �����  �  H         ����
    !           u � 6f       �����F  �      l     �� ��^       ����	 � �����  �  H         ����
  " #           y � =j       �����G  ��      l     �� ��^       ����	 � �����  �  H         ����
  $ %           } � Dn       �����H  ,�      l     �� ��^       ����	 � �����  �  H         ����
  & '           � � Kr       �����I  ��      l     �� ��^       ����	 � �����  �  H         ����
  ( )           � � Rv       �����J  D�      l     �� ��^       ����	 � �����  �  H         ����
  * +           � � Yz       �����K  ��       l     �� ��^       ����	 � �����  �  H         ����
  , -           � � `~       �����L  \    ��  l	     �� ��^       ����	 � �����  �  H          ����              " % . (       �����  X       �      �� ��_        ���� � ������������I          ����              $ ( 3 *       ����  $       �     �� ��_        ���� � ������������I          ����              & + 8 ,       ����0  `       �     �� ��_        ���� � ������������I          ����   	           ( . = .       ����N  �       �     �� ��_       ���� � ������������I          ����  
            * 1 B 0       ����l  �       �     �� ��_       ���� � ������������I          ����              , 4 G 2       �����         �     �� ��_       ���� � ������������I          ����              . 7 L 4       �����  P       �     �� ��_       ���� � ������������I          ����              0 : Q 6       �����  �       �     �� ��_       ���� � ������������I          ����              2 = V 8       �����  �       �     �� ��_       ���� � ������������I          ����              4 @ [ :       ����         �	     �� ��_       ���� � ������������I          ����              & - I +       ����z  n
       �      �� ��`        ���� � ������������J          ����              ) 0 N -       �����  "       �     �� ��`        ���� � ������������J          ����  	 
           , 3 S /       �����  �       �     �� ��`        ���� � ������������J          ����              / 6 X 1       ����.  �       �     �� ��`       ���� � ������������J          ����              2 9 ] 3       ����j  >       �     �� ��`       ���� � ������������J          ����              5 < b 5       �����  �       �     �� ��`       ���� � ������������J          ����              8 ? g 7       �����  �       �     �� ��`       ���� � ������������J          ����              ; B l 9       ����  Z       �     �� ��`       ���� � ������������J          ����              > E q ;       ����Z         �     �� ��`       ���� � ������������J          ����              A H v =       �����  �       �	     �� ��`       ���� � ������������J         ����   	           * 4 c .       �����         �      �� ��a        ���� � ������������K         ����  
            - 8 h 1       �����  �       �     �� ��a        ���� � ������������K         ����              0 < m 4       ����:  �       �     �� ��a        ���� � ������������K         ����              3 @ r 7       �����  P       �     �� ��a       ���� � ������������K         ����              6 D w :       �����  �       �     �� ��a       ���� � ������������K         ����              9 H | =       ����H   !       �     �� ��a       ���� � ������������K         ����              < L � @       �����  �"       �     �� ��a       ���� � ������������K         ����              ? P � C       �����  �#       �     �� ��a       ���� � ������������K         ����              B T � F       ����V	  X%       �     �� ��a       ���� � ������������K         ����              E X � I       �����	  �&       �	     �� ��a       ���� � ������������K         ����              2 E | 6       ����  x7       �      �� ��b        ���� � ������������L         ����              5 I � 9       �����  �9       �     �� ��b        ���� � ������������L         ����              8 M � <       ����  (<       �     �� ��b        ���� � ������������L         ����              ; Q � ?       �����  �>       �     �� ��b       ���� � ������������L         ����              > U � B       �����  �@       �     �� ��b       ���� � ������������L         ����              A Y � E       ����p  0C       �     �� ��b       ���� � ������������L         ����              D ] � H       �����  �E       �     �� ��b       ���� � ������������L         ����              G a � K       ����`  �G       �     �� ��b       ���� � ������������L         ����              J e � N       �����  8J       �     �� ��b       ���� � ������������L         ����              M i � Q       ����P  �L       �	     �� ��b       ���� � ������������L         ����              9 U � =       ����0   g       �      �� ��c        ���� � ������������M         ����              < Y � @       �����  �j       �     �� ��c        ���� � ������������M         ����              ? ] � C       ����\  (n       �     �� ��c        ���� � ������������M         ����              B a � F       �����  �q       �     �� ��c       ���� � ������������M         ����              E e � I       �����  0u       �     �� ��c       ���� � ������������M         ����              H i � L       ����  �x       �     �� ��c       ���� � ������������M         ����              K m � O       �����  8|       �     �� ��c       ���� � ������������M         ����              N q � R       ����J  �       �     �� ��c       ���� � ������������M         ����              Q u � U       �����  @�    
   �     �� ��c       ���� � ������������M         ����    !           T y � X       ����v  Ć    	   �	     �� ��c       ���� � ������������M         ����              @ d � D       �����  ��       �      �� ��d        ���� � ������������N         ����              D h � G       �����  ��       �     �� ��d        ���� � ������������N         ����              H l � J       ����6  z�       �     �� ��d        ���� � ������������N         ����              L p � M       �����  f�       �     �� ��d       ���� � ������������N         ����              P t � P       �����  R�       �     �� ��d       ���� � ������������N         ����              T x � S       ����R  >�       �     �� ��d       ���� � ������������N         ����              X | � V       ����  *�       �     �� ��d       ���� � ������������N         ����               \ � � Y       �����  �    	   �     �� ��d       ���� � ������������N         ����  ! "           ` � � \       ����n  �       �     �� ��d       ���� � ������������N         ����  # $           d � � _       ����"  ��       �	     �� ��d       ���� � ������������N         ����              P s � J       �����!  �      �      �� ��e        ���� � �����  �  O         ����              T x � N       �����"         �     �� ��e        ���� � �����  �  O         ����              X } � R       �����#  �      �     �� ��e        ���� � �����  �  O         ����              \ � � V       ����h$  @#      �     �� ��e       ���� � �����  �  O         ����              ` � � Z       ����:%  �)      �     �� ��e       ���� � �����  �  O         ����              d � � ^       ����&  `0   	   �     �� ��e       ���� � �����  �  O         ����    !           h � b       �����&  �6      �     �� ��e       ���� � �����  �  O         ����  " #           l � f       �����'  �=      �     �� ��e       ���� � �����  �  O         ����  $ %           p � j       �����(  D      �     �� ��e       ���� � �����  �  O         ����  & '           t � n       ����T)  �J      �	     �� ��e       ���� � �����  �  O         ����              ` � Z       �����,  |�      �      �� ��f        ���� � �����  �  P         ����              d � ^       �����-  �      �     �� ��f        ���� � �����  �  P         ����              h � b       ����|.  \�      �     �� ��f        ���� � �����  �  P         ����              l � f       ����l/  ̪   	   �     �� ��f       ���� � �����  �  P         ����               p � j       ����\0  <�      �     �� ��f       ���� � �����  �  P         ����  ! "           t � $n       ����L1  ��      �     �� ��f       ���� � �����  �  P         ����  # $           x � +r       ����<2  �      �     �� ��f       ���� � �����  �  P         ����  % &           | � 2v       ����,3  ��      �     �� ��f       ���� � �����  �  P         ����  ' (           � � 9z       ����4  ��      �     �� ��f       ���� � �����  �  P         ����  ) *           � � @~       ����5  l�      �	     �� ��f       ���� � �����  �  P         ����              o � *i       �����8  �7      �      �� ��g        ����	 � �����  �  Q         ����              s � 1m       �����9  �B   
   �     �� ��g        ����	 � �����  �  Q         ����              w � 8q       �����:  M      �     �� ��g        ����	 � �����  �  Q         ����    !           { � ?u       �����;  �W      �     �� ��g       ����	 � �����  �  Q         ����  " #            � Fy       ����=  (b      �     �� ��g       ����	 � �����  �  Q         ����  $ %           � � M}       ����>  �l      �     �� ��g       ����	 � �����  �  Q         ����  & '           � � T�       ���� ?  @w      �     �� ��g       ����	 � �����  �  Q         ����  ( )           � � [�       ����.@  ́      �     �� ��g       ����	 � �����  �  Q         ����  * +           � � b�       ����<A  X�       �     �� ��g       ����	 � �����  �  Q         ����  , -           � � i�       ����JB  �   ��  �	     �� ��g       ����	 � �����  �  Q          ����              + . 7 1       �����  �              �� ��h        ���� � ������������R          ����              - 1 < 3       �����  |            �� ��h        ���� � ������������R          ����              / 4 A 5       �����  �            �� ��h        ���� � ������������R          ����   	           1 7 F 7       �����  �            �� ��h       ���� � ������������R          ����  
            3 : K 9       ����  0             �� ��h       ���� � ������������R          ����              5 = P ;       ����6  l             �� ��h       ���� � ������������R          ����              7 @ U =       ����T  �             �� ��h       ���� � ������������R          ����              9 C Z ?       ����r  �             �� ��h       ���� � ������������R          ����              ; F _ A       �����   !            �� ��h       ���� � ������������R          ����              = I d C       �����  \!       	     �� ��h       ���� � ������������R          ����              - 6 R 3       ����&  r3             �� ��i        ���� � ������������S          ����              0 9 W 5       ����b  &4            �� ��i        ���� � ������������S          ����  	 
           3 < \ 7       �����  �4            �� ��i        ���� � ������������S          ����              6 ? a 9       �����  �5            �� ��i       ���� � ������������S          ����              9 B f ;       ����  B6            �� ��i       ���� � ������������S          ����              < E k =       ����R  �6            �� ��i       ���� � ������������S          ����              ? H p ?       �����  �7            �� ��i       ���� � ������������S          ����              B K u A       �����  ^8            �� ��i       ���� � ������������S          ����              E N z C       ����  9            �� ��i       ���� � ������������S          ����              H Q  E       ����B  �9       	     �� ��i       ���� � ������������S         ����   	           / = l 5       ����2  �P             �� ��j        ���� � ������������T         ����  
            2 A q 8       �����  0R            �� ��j        ���� � ������������T         ����              5 E v ;       �����  �S            �� ��j        ���� � ������������T         ����              8 I { >       ����@   U            �� ��j       ���� � ������������T         ����              ; M � A       �����  hV            �� ��j       ���� � ������������T         ����              > Q � D       �����  �W            �� ��j       ���� � ������������T         ����              A U � G       ����N  8Y            �� ��j       ���� � ������������T         ����              D Y � J       �����  �Z            �� ��j       ���� � ������������T         ����              G ] � M       ����  \            �� ��j       ���� � ������������T         ����              J a � P       ����\  p]       	     �� ��j       ���� � ������������T         ����              7 N � 7       �����  �{             �� ��k        ���� � ������������U         ����              : R � :       ����<  ,~            �� ��k        ���� � ������������U         ����              = V � =       �����  ��            �� ��k        ���� � ������������U         ����              @ Z � @       ����,  ܂            �� ��k       ���� � ������������U         ����              C ^ � C       �����  4�            �� ��k       ���� � ������������U         ����              F b � F       ����  ��            �� ��k       ���� � ������������U         ����              I f � I       �����  �            �� ��k       ���� � ������������U         ����              L j � L       ����  <�            �� ��k       ���� � ������������U         ����              O n � O       �����  ��            �� ��k       ���� � ������������U         ����              R r � R       �����  �       	     �� ��k       ���� � ������������U         ����              > ^ � >       �����  (�             �� ��l        ���� � ������������V         ����              A b � A       ����r  ��            �� ��l        ���� � ������������V         ����              D f � D       ����   0�            �� ��l        ���� � ������������V         ����              G j � G       �����   ��            �� ��l       ���� � ������������V         ����              J n � J       ����4!  8�            �� ��l       ���� � ������������V         ����              M r � M       �����!  ��            �� ��l       ���� � ������������V         ����              P v � P       ����`"  @�            �� ��l       ���� � ������������V         ����              S z � S       �����"  ��            �� ��l       ���� � ������������V         ����              V ~ � V       �����#  H�    
        �� ��l       ���� � ������������V         ����    !           Y � � Y       ����"$  ��    	   	     �� ��l       ���� � ������������V         ����              E m � E       ����z&  V            �� ��m        ���� � ������������W         ����              I q � H       ����.'  B           �� ��m        ���� � ������������W         ����              M u � K       �����'  .           �� ��m        ���� � ������������W         ����              Q y � N       �����(             �� ��m       ���� � ������������W         ����              U } � Q       ����J)  !           �� ��m       ���� � ������������W         ����              Y � � T       �����)  �%           �� ��m       ���� � ������������W         ����              ] � � W       �����*  �*           �� ��m       ���� � ������������W         ����               a � � Z       ����f+  �/   	        �� ��m       ���� � ������������W         ����  ! "           e � � ]       ����,  �4           �� ��m       ���� � ������������W         ����  # $           i � � `       �����,  �9      	     �� ��m       ���� � ������������W         ����              U | � K       �����/  �|            �� ��n        ���� � �����  �  X         ����              Y � � O       ����p0  ��           �� ��n        ���� � �����  �  X         ����              ] � � S       ����B1  �           �� ��n        ���� � �����  �  X         ����              a � � W       ����2  ��           �� ��n       ���� � �����  �  X         ����              e � [       �����2  0�           �� ��n       ���� � �����  �  X         ����              i � _       �����3  ��   	        �� ��n       ���� � �����  �  X         ����    !           m � c       �����4  P�           �� ��n       ���� � �����  �  X         ����  " #           q � g       ����\5  �           �� ��n       ���� � �����  �  X         ����  $ %           u � k       ����.6  p�           �� ��n       ���� � �����  �  X         ����  & '           y �  o       ���� 7   �      	     �� ��n       ���� � �����  �  X         ����              e � 
[       ����H:  �            �� ��o        ���� � �����  �  Y         ����              i � _       ����8;  �           �� ��o        ���� � �����  �  Y         ����              m � c       ����(<  h           �� ��o        ���� � �����  �  Y         ����              q � g       ����=  �%   	        �� ��o       ���� � �����  �  Y         ����               u � &k       ����>  H.           �� ��o       ���� � �����  �  Y         ����  ! "           y � -o       �����>  �6           �� ��o       ���� � �����  �  Y         ����  # $           } � 4s       �����?  (?           �� ��o       ���� � �����  �  Y         ����  % &           � � ;w       �����@  �G           �� ��o       ���� � �����  �  Y         ����  ' (           � � B{       �����A  P           �� ��o       ���� � �����  �  Y         ����  ) *           � � I       �����B  xX      	     �� ��o       ���� � �����  �  Y         ����              t � 3j       ����xF  ��             �� ��p        ����	 � �����  �  Z         ����              x � :n       �����G  <�   
         �� ��p        ����	 � �����  �  Z         ����              | � Ar       �����H  ��            �� ��p        ����	 � �����  �  Z         ����    !           � � Hv       �����I  T�            �� ��p       ����	 � �����  �  Z         ����  " #           � � Oz       �����J  ��            �� ��p       ����	 � �����  �  Z         ����  $ %           � � V~       �����K  l�            �� ��p       ����	 � �����  �  Z         ����  & '           � � ]�       �����L  ��            �� ��p       ����	 � �����  �  Z         ����  ( )           � � d�       �����M  �
            �� ��p       ����	 � �����  �  Z         ����  * +           � � k�       �����N               �� ��p       ����	 � �����  �  Z         ����  , -           � � r�       �����O  �   ��   	     �� ��p       ����	 � �����  �  Z          ����              . 1 : 4       ����0  �        r      �� ��q        ���� � ������������[          ����              0 4 ? 6       ����N  �"       r     �� ��q        ���� � ������������[          ����              2 7 D 8       ����l  �"       r     �� ��q        ���� � ������������[          ����   	           4 : I :       �����  #       r     �� ��q       ���� � ������������[          ����  
            6 = N <       �����  P#       r     �� ��q       ���� � ������������[          ����              8 @ S >       �����  �#       r     �� ��q       ���� � ������������[          ����              : C X @       �����  �#       r     �� ��q       ���� � ������������[          ����              < F ] B       ����  $       r     �� ��q       ���� � ������������[          ����              > I b D       ����   @$       r     �� ��q       ���� � ������������[          ����              @ L g F       ����>  |$       r	     �� ��q       ���� � ������������[          ����              1 9 U 6       �����  "8       s      �� ��r        ���� � ������������\          ����              4 < Z 8       �����  �8       s     �� ��r        ���� � ������������\          ����  	 
           7 ? _ :       ����.  �9       s     �� ��r        ���� � ������������\          ����              : B d <       ����j  >:       s     �� ��r       ���� � ������������\          ����              = E i >       �����  �:       s     �� ��r       ���� � ������������\          ����              @ H n @       �����  �;       s     �� ��r       ���� � ������������\          ����              C K s B       ����  Z<       s     �� ��r       ���� � ������������\          ����              F N x D       ����Z  =       s     �� ��r       ���� � ������������\          ����              I Q } F       �����  �=       s     �� ��r       ���� � ������������\          ����              L T � H       �����  v>       s	     �� ��r       ���� � ������������\         ����   	           9 @ o 8       �����  W       t      �� ��s        ���� � ������������]         ����  
            < D t ;       ����  pX       t     �� ��s        ���� � ������������]         ����              ? H y >       ����v  �Y       t     �� ��s        ���� � ������������]         ����              B L ~ A       �����  @[       t     �� ��s       ���� � ������������]         ����              E P � D       ����*  �\       t     �� ��s       ���� � ������������]         ����              H T � G       �����  ^       t     �� ��s       ���� � ������������]         ����              K X � J       �����  x_       t     �� ��s       ���� � ������������]         ����              N \ � M       ����8  �`       t     �� ��s       ���� � ������������]         ����              Q ` � P       �����  Hb       t     �� ��s       ���� � ������������]         ����              T d � S       �����  �c       t	     �� ��s       ���� � ������������]         ����              A Q � <       ����T  ��       u      �� ��t        ���� � ������������^         ����              D U � ?       �����  ��       u     �� ��t        ���� � ������������^         ����              G Y � B       ����D  T�       u     �� ��t        ���� � ������������^         ����              J ] � E       �����  ��       u     �� ��t       ���� � ������������^         ����              M a � H       ����4  �       u     �� ��t       ���� � ������������^         ����              P e � K       �����  \�       u     �� ��t       ���� � ������������^         ����              S i � N       ����$  ��       u     �� ��t       ���� � ������������^         ����              V m � Q       �����  �       u     �� ��t       ���� � ������������^         ����              Y q � T       ����  d�       u     �� ��t       ���� � ������������^         ����              \ u � W       �����  ��       u	     �� ��t       ���� � ������������^         ����              H a � C       ����l   ��       v      �� ��u        ���� � ������������_         ����              K e � F       ����!  �       v     �� ��u        ���� � ������������_         ����              N i � I       �����!  ��       v     �� ��u        ���� � ������������_         ����              Q m � L       ����."  �       v     �� ��u       ���� � ������������_         ����              T q � O       �����"  ��       v     �� ��u       ���� � ������������_         ����              W u � R       ����Z#  �       v     �� ��u       ���� � ������������_         ����              Z y � U       �����#  ��       v     �� ��u       ���� � ������������_         ����              ] } � X       �����$  $�       v     �� ��u       ���� � ������������_         ����              ` � � [       ����%  ��    
   v     �� ��u       ���� � ������������_         ����    !           c � � ^       �����%  ,�    	   v	     �� ��u       ���� � ������������_         ����              O p � J       ����
(  F      w      �� ��v        ���� � ������������`         ����              S t � M       �����(  2      w     �� ��v        ���� � ������������`         ����              W x � P       ����r)  "      w     �� ��v        ���� � ������������`         ����              [ | � S       ����&*  
'      w     �� ��v       ���� � ������������`         ����              _ � � V       �����*  �+      w     �� ��v       ���� � ������������`         ����              c � � Y       �����+  �0      w     �� ��v       ���� � ������������`         ����              g � � \       ����B,  �5      w     �� ��v       ���� � ������������`         ����               k � � _       �����,  �:   	   w     �� ��v       ���� � ������������`         ����  ! "           o � � b       �����-  �?      w     �� ��v       ���� � ������������`         ����  # $           s � e       ����^.  �D      w	     �� ��v       ���� � ������������`         ����              _  � P       ����.1  p�      x      �� ��w        ���� � �����  �  a         ����              c � � T       ���� 2   �      x     �� ��w        ���� � �����  �  a         ����              g � � X       �����2  ��      x     �� ��w        ���� � �����  �  a         ����              k � � \       �����3   �      x     �� ��w       ���� � �����  �  a         ����              o � `       ����v4  ��      x     �� ��w       ���� � �����  �  a         ����              s � d       ����H5  @�   	   x     �� ��w       ���� � �����  �  a         ����    !           w � h       ����6  а      x     �� ��w       ���� � �����  �  a         ����  " #           { � l       �����6  `�      x     �� ��w       ���� � �����  �  a         ����  $ %            � p       �����7  �      x     �� ��w       ���� � �����  �  a         ����  & '           � � #t       �����8  ��      x	     �� ��w       ���� � �����  �  a         ����              o � `       �����;  �      y      �� ��x        ���� � �����  �  b         ����              s � d       �����<  #      y     �� ��x        ���� � �����  �  b         ����              w � h       �����=  x+      y     �� ��x        ���� � �����  �  b         ����              { � "l       �����>  �3   	   y     �� ��x       ���� � �����  �  b         ����                � )p       �����?  X<      y     �� ��x       ���� � �����  �  b         ����  ! "           � � 0t       �����@  �D      y     �� ��x       ���� � �����  �  b         ����  # $           � � 7x       ����xA  8M      y     �� ��x       ���� � �����  �  b         ����  % &           � � >|       ����hB  �U      y     �� ��x       ���� � �����  �  b         ����  ' (           � � E�       ����XC  ^      y     �� ��x       ���� � �����  �  b         ����  ) *           � � L�       ����HD  �f      y	     �� ��x       ���� � �����  �  b         ����              ~ � 6o       ����H  P�      z      �� ��y        ����	 � �����  �  c         ����              � � =s       ����I  ��   
   z     �� ��y        ����	 � �����  �  c         ����              � � Dw       ����$J  h�      z     �� ��y        ����	 � �����  �  c         ����    !           � � K{       ����2K  ��      z     �� ��y       ����	 � �����  �  c         ����  " #           � � R       ����@L  ��      z     �� ��y       ����	 � �����  �  c         ����  $ %           � � Y�       ����NM        z     �� ��y       ����	 � �����  �  c         ����  & '           � � `�       ����\N  �      z     �� ��y       ����	 � �����  �  c         ����  ( )           � � g�       ����jO  $      z     �� ��y       ����	 � �����  �  c         ����  * +           � � n�       ����xP  �$       z     �� ��y       ����	 � �����  �  c         ����  , -           � � u�       �����Q  </   ��  z	     �� ��y       ����	 � �����  �  c          ��  3 4           l� h \ x     ����~O  jj       �       �    z        ����
 � �����  �  d          ��  5 6           s� l ` x     �����P  Nw       �      �    z        ����
 � �����  �  d          ��  7 8           z� p d x     �����Q  2�       �      �    z        ����
 � �����  �  d          ��  : ;           �� t h x     ����S  �       �      �    z        ����
 � �����  �  d          ��  < =           �� x l x     ����.T  ��       �      �    z        ����
 � �����  �  d          ��  > ?           �� | p x     ����ZU  ު       �      �    z        ����
 � �����  �  d          ��  @ A           �� � t x     �����V  ·       �      �    z        ����
 � �����  �  d          ��  B C           �� � x x     �����W  ��       �      �    z        ����
 � �����  �  d          ��  E F           �� � | x     �����X  ��       �      �    z        ����
 � �����  �  d          ��  G H           �� � � x     ����
Z  n�       � 	     �    z        ����
 �����  �  d          ��  ' (           � � eb x     ����~O  jj       �       �    {        ����
 � �����  �  e          ��  ) *           � � lf x     �����P  Nw       �      �    {        ����
 � �����  �  e          ��  + ,           � � sj x     �����Q  2�       �      �    {        ����
 � �����  �  e          ��  - .           � � zn x     ����S  �       �      �    {        ����
 � �����  �  e          ��  / 0           � � �r x     ����.T  ��       �      �    {        ����
 � �����  �  e          ��  1 2           � � �v x     ����ZU  ު       �      �    {        ����
 � �����  �  e          ��  4 5           � � �z x     �����V  ·       �      �    {        ����
 � �����  �  e          ��  6 7           � � �~ x     �����W  ��       �      �    {        ����
 � �����  �  e          ��  8 9           � � �� x     �����X  ��       �      �    {        ����
 � �����  �  e          ��  : ;           � �� x     ����
Z  n�       � 	     �    {        ����
 �����  �  e          ��  & '           ([ (] x     ����~O  jj       �       �    |        ����
 � �����  �  f          ��  ( )           ._ .a x     �����P  Nw       �      �    |        ����
 � �����  �  f          ��  * +           4c 4e x     �����Q  2�       �      �    |        ����
 � �����  �  f          ��  , -           :g :i x     ����S  �       �      �    |        ����
 � �����  �  f          ��  . /           @k @m x     ����.T  ��       �      �    |        ����
 � �����  �  f          ��  0 1           Fo Fq x     ����ZU  ު       �      �    |        ����
 � �����  �  f          ��  3 4           Ls Lu x     �����V  ·       �      �    |        ����
 � �����  �  f          ��  5 6           Rw Ry x     �����W  ��       �      �    |        ����
 � �����  �  f          ��  7 8           X{ X} x     �����X  ��       �      �    |        ����
 � �����  �  f          ��  9 :           ^ ^� x     ����
Z  n�       � 	     �    |        ����
 �����  �  f          ��              � � Xv x     ����~O  jj       �       �    }        ����
 � �����  �  g          ��               � � _z x     �����P  Nw       �      �    }        ����
 � �����  �  g          ��  ! "           � � f~ x     �����Q  2�       �      �    }        ����
 � �����  �  g          ��  # $           � � m� x     ����S  �       �      �    }        ����
 � �����  �  g          ��  % &           � � t� x     ����.T  ��       �      �    }        ����
 � �����  �  g          ��  ' (           � � {� x     ����ZU  ު       �      �    }        ����
 � �����  �  g          ��  ) *           � � �� x     �����V  ·       �      �    }        ����
 � �����  �  g          ��  + ,           � � �� x     �����W  ��       �      �    }        ����
 � �����  �  g          ��  - .           � � �� x     �����X  ��       �      �    }        ����
 � �����  �  g          ��  / 0           � � �� x     ����
Z  n�       � 	     �    }        ����
 �����  �  g         ����	  0 1           H� h \       �����R  ʌ   	   �      �� ��~        ����
 � �����  �  h         ����	  2 3           O� l `       �����S  ��      �     �� ��~        ����
 � �����  �  h         ����	  4 5           V� p d       �����T  ��      �     �� ��~        ����
 � �����  �  h         ����	  7 8           ]� t h       ����"V  v�      �     �� ��~       ����
 � �����  �  h         ����	  9 :           d� x l       ����NW  Z�      �     �� ��~       ����
 � �����  �  h         ����	  ; <           k� | p       ����zX  >�      �     �� ��~       ����
 � �����  �  h         ����	  = >           r� � t       �����Y  "�      �     �� ��~       ����
 � �����  �  h         ����	  ? @           y� � x       �����Z  �   ��  �     �� ��~       ����
 � �����  �  h         ����	  B C           �� � |       �����[  ��   ��  �     �� ��~       ����
 � �����  �  h         ����	  D E           �� � �       ����*]  �    ��  �	     �� ��~       ����
 �����  �  h         ����	  & '           t � Ab       �����R  ʌ   	   �      �� ��        ����
 � �����  �  i         ����	  ( )           y � Hf       �����S  ��      �     �� ��        ����
 � �����  �  i         ����	  * +           ~ � Oj       �����T  ��      �     �� ��        ����
 � �����  �  i         ����	  , -           � � Vn       ����"V  v�      �     �� ��       ����
 � �����  �  i         ����	  . /           � � ]r       ����NW  Z�      �     �� ��       ����
 � �����  �  i         ����	  0 1           � � dv       ����zX  >�      �     �� ��       ����
 � �����  �  i         ����	  3 4           � � kz       �����Y  "�      �     �� ��       ����
 � �����  �  i         ����	  5 6           � � r~       �����Z  �   ��  �     �� ��       ����
 � �����  �  i         ����	  7 8           � � y�       �����[  ��   ��  �     �� ��       ����
 � �����  �  i         ����	  9 :           � � ��       ����*]  �    ��  �	     �� ��       ����
 �����  �  i         ����	  % &           [ ]       �����R  ʌ   	         �� ���        ����
 � �����  �  j         ����	  ' (           
_ 
a       �����S  ��           �� ���        ����
 � �����  �  j         ����	  ) *           c e       �����T  ��           �� ���        ����
 � �����  �  j         ����	  + ,           g i       ����"V  v�           �� ���       ����
 � �����  �  j         ����	  - .           k m       ����NW  Z�           �� ���       ����
 � �����  �  j         ����	  / 0           "o "q       ����zX  >�           �� ���       ����
 � �����  �  j         ����	  2 3           (s (u       �����Y  "�           �� ���       ����
 � �����  �  j         ����	  4 5           .w .y       �����Z  �   ��       �� ���       ����
 � �����  �  j         ����	  6 7           4{ 4}       �����[  ��   ��       �� ���       ����
 � �����  �  j         ����	  8 9           : :�       ����*]  �    ��  	     �� ���       ����
 �����  �  j         ����	              q � @`       �����R  ʌ   	         �� ���        ����
 � �����  �  k         ����	               v � Gd       �����S  ��           �� ���        ����
 � �����  �  k         ����	  ! "           { � Nh       �����T  ��           �� ���        ����
 � �����  �  k         ����	  # $           � � Ul       ����"V  v�           �� ���       ����
 � �����  �  k         ����	  % &           � � \p       ����NW  Z�           �� ���       ����
 � �����  �  k         ����	  ' (           � � ct       ����zX  >�           �� ���       ����
 � �����  �  k         ����	  ) *           � � jx       �����Y  "�           �� ���       ����
 � �����  �  k         ����	  + ,           � � q|       �����Z  �   ��       �� ���       ����
 � �����  �  k         ����	  - .           � � x�       �����[  ��   ��       �� ���       ����
 � �����  �  k         ����	  / 0           � � �       ����*]  �    ��  	     �� ���       ����
 �����  �  k         ����
  1 2           U� h \       ����Q  �{   	   @      �� ���        ����
 � �����  �  l         ����
  3 4           \� l `       ����:R  ~�      @     �� ���        ����
 � �����  �  l         ����
  5 6           c� p d       ����fS  b�      @     �� ���        ����
 � �����  �  l         ����
  8 9           j� t h       �����T  F�      @     �� ���       ����
 � �����  �  l         ����
  : ;           q� x l       �����U  *�      @     �� ���       ����
 � �����  �  l         ����
  < =           x� | p       �����V  �      @     �� ���       ����
 � �����  �  l         ����
  > ?           � � t       ����X  ��      @     �� ���       ����
 � �����  �  l         ����
  @ A           �� � x       ����BY  ��   ��  @     �� ���       ����
 � �����  �  l         ����
  C D           �� � |       ����nZ  ��   ��  @     �� ���       ����
 � �����  �  l         ����
  E F           �� � �       �����[  ��   ��  @	     �� ���       ����
 �����  �  l         ����
  & '           � � Nb       ����Q  �{   	   O      �� ���        ����
 � �����  �  m         ����
  ( )           � � Uf       ����:R  ~�      O     �� ���        ����
 � �����  �  m         ����
  * +           � � \j       ����fS  b�      O     �� ���        ����
 � �����  �  m         ����
  , -           � � cn       �����T  F�      O     �� ���       ����
 � �����  �  m         ����
  . /           � � jr       �����U  *�      O     �� ���       ����
 � �����  �  m         ����
  0 1           � � qv       �����V  �      O     �� ���       ����
 � �����  �  m         ����
  3 4           � � xz       ����X  ��      O     �� ���       ����
 � �����  �  m         ����
  5 6           � � ~       ����BY  ��   ��  O     �� ���       ����
 � �����  �  m         ����
  7 8           � � ��       ����nZ  ��   ��  O     �� ���       ����
 � �����  �  m         ����
  9 :           � � ��       �����[  ��   ��  O	     �� ���       ����
 �����  �  m         ����
  % &           [ ]       ����Q  �{   	   ^      �� ���        ����
 � �����  �  n         ����
  ' (           _ a       ����:R  ~�      ^     �� ���        ����
 � �����  �  n         ����
  ) *           c e       ����fS  b�      ^     �� ���        ����
 � �����  �  n         ����
  + ,           #g #i       �����T  F�      ^     �� ���       ����
 � �����  �  n         ����
  - .           )k )m       �����U  *�      ^     �� ���       ����
 � �����  �  n         ����
  / 0           /o /q       �����V  �      ^     �� ���       ����
 � �����  �  n         ����
  2 3           5s 5u       ����X  ��      ^     �� ���       ����
 � �����  �  n         ����
  4 5           ;w ;y       ����BY  ��   ��  ^     �� ���       ����
 � �����  �  n         ����
  6 7           A{ A}       ����nZ  ��   ��  ^     �� ���       ����
 � �����  �  n         ����
  8 9           G G�       �����[  ��   ��  ^	     �� ���       ����
 �����  �  n         ����
              x � Ii       ����Q  �{   	   m      �� ���        ����
 � �����  �  o         ����
               } � Pm       ����:R  ~�      m     �� ���        ����
 � �����  �  o         ����
  ! "           � � Wq       ����fS  b�      m     �� ���        ����
 � �����  �  o         ����
  # $           � � ^u       �����T  F�      m     �� ���       ����
 � �����  �  o         ����
  % &           � � ey       �����U  *�      m     �� ���       ����
 � �����  �  o         ����
  ' (           � � l}       �����V  �      m     �� ���       ����
 � �����  �  o         ����
  ) *           � � s�       ����X  ��      m     �� ���       ����
 � �����  �  o         ����
  + ,           � � z�       ����BY  ��   ��  m     �� ���       ����
 � �����  �  o         ����
  - .           � � ��       ����nZ  ��   ��  m     �� ���       ����
 � �����  �  o         ����
  / 0           � � ��       �����[  ��   ��  m	     �� ���       ����
 �����  �  o         ����  2 3           b� h \       �����F  �   	   �      �� ���        ����
 � �����  �  p         ����  4 5           i� l `       �����G  z      �     �� ���        ����
 � �����  �  p         ����  6 7           p� p d       �����H  ^!      �     �� ���        ����
 � �����  �  p         ����  9 :           w� t h       ����J  B.      �     �� ���       ����
 � �����  �  p         ����  ; <           ~� x l       ����2K  &;      �     �� ���       ����
 � �����  �  p         ����  = >           �� | p       ����^L  
H      �     �� ���       ����
 � �����  �  p         ����  ? @           �� � t       �����M  �T      �     �� ���       ����
 � �����  �  p         ����  A B           �� � x       �����N  �a   ��  �     �� ���       ����
 � �����  �  p         ����  D E           �� � |       �����O  �n   ��  �     �� ���       ����
 � �����  �  p         ����  F G           �� � �       ����Q  �{   ��  �	     �� ���       ����
 �����  �  p         ����  ' (           � � [b       �����F  �   	   �      �� ���        ����
 � �����  �  q         ����  ) *           � � bf       �����G  z      �     �� ���        ����
 � �����  �  q         ����  + ,           � � ij       �����H  ^!      �     �� ���        ����
 � �����  �  q         ����  - .           � � pn       ����J  B.      �     �� ���       ����
 � �����  �  q         ����  / 0           � � wr       ����2K  &;      �     �� ���       ����
 � �����  �  q         ����  1 2           � � ~v       ����^L  
H      �     �� ���       ����
 � �����  �  q         ����  4 5           � � �z       �����M  �T      �     �� ���       ����
 � �����  �  q         ����  6 7           � � �~       �����N  �a   ��  �     �� ���       ����
 � �����  �  q         ����  8 9           � � ��       �����O  �n   ��  �     �� ���       ����
 � �����  �  q         ����  : ;           � � ��       ����Q  �{   ��  �	     �� ���       ����
 �����  �  q         ����  & '           [ ]       �����F  �   	   �      �� ���        ����
 � �����  �  r         ����  ( )           $_ $a       �����G  z      �     �� ���        ����
 � �����  �  r         ����  * +           *c *e       �����H  ^!      �     �� ���        ����
 � �����  �  r         ����  , -           0g 0i       ����J  B.      �     �� ���       ����
 � �����  �  r         ����  . /           6k 6m       ����2K  &;      �     �� ���       ����
 � �����  �  r         ����  0 1           <o <q       ����^L  
H      �     �� ���       ����
 � �����  �  r         ����  3 4           Bs Bu       �����M  �T      �     �� ���       ����
 � �����  �  r         ����  5 6           Hw Hy       �����N  �a   ��  �     �� ���       ����
 � �����  �  r         ����  7 8           N{ N}       �����O  �n   ��  �     �� ���       ����
 � �����  �  r         ����  9 :           T T�       ����Q  �{   ��  �	     �� ���       ����
 �����  �  r         ����              ~ � Rx       �����F  �   	   �      �� ���        ����
 � �����  �  s         ����               � � Y|       �����G  z      �     �� ���        ����
 � �����  �  s         ����  ! "           � � `�       �����H  ^!      �     �� ���        ����
 � �����  �  s         ����  # $           � � g�       ����J  B.      �     �� ���       ����
 � �����  �  s         ����  % &           � � n�       ����2K  &;      �     �� ���       ����
 � �����  �  s         ����  ' (           � � u�       ����^L  
H      �     �� ���       ����
 � �����  �  s         ����  ) *           � � |�       �����M  �T      �     �� ���       ����
 � �����  �  s         ����  + ,           � � ��       �����N  �a   ��  �     �� ���       ����
 � �����  �  s         ����  - .           � � ��       �����O  �n   ��  �     �� ���       ����
 � �����  �  s         ����  / 0           � � ��       ����Q  �{   ��  �	     �� ���       ����
 �����  �  s         ����  3 4           o� h \       ����.T  ��   	   �      �� ���        ����
 � �����  �  t         ����  5 6           v� l `       ����ZU  ު      �     �� ���        ����
 � �����  �  t         ����  7 8           }� p d       �����V  ·      �     �� ���        ����
 � �����  �  t         ����  : ;           �� t h       �����W  ��      �     �� ���       ����
 � �����  �  t         ����  < =           �� x l       �����X  ��      �     �� ���       ����
 � �����  �  t         ����  > ?           �� | p       ����
Z  n�      �     �� ���       ����
 � �����  �  t         ����  @ A           �� � t       ����6[  R�      �     �� ���       ����
 � �����  �  t         ����  B C           �� � x       ����b\  6�   ��  �     �� ���       ����
 � �����  �  t         ����  E F           �� � |       �����]     ��  �     �� ���       ����
 � �����  �  t         ����  G H           �� � �       �����^  �   ��  �	     �� ���       ����
 �����  �  t         ����  ' (           � � hb       ����.T  ��   	         �� ���        ����
 � �����  �  u         ����  ) *           � � of       ����ZU  ު           �� ���        ����
 � �����  �  u         ����  + ,           � � vj       �����V  ·           �� ���        ����
 � �����  �  u         ����  - .           � � }n       �����W  ��           �� ���       ����
 � �����  �  u         ����  / 0           � � �r       �����X  ��           �� ���       ����
 � �����  �  u         ����  1 2           � � �v       ����
Z  n�           �� ���       ����
 � �����  �  u         ����  4 5           � � �z       ����6[  R�           �� ���       ����
 � �����  �  u         ����  6 7           � � �~       ����b\  6�   ��       �� ���       ����
 � �����  �  u         ����  8 9           � � ��       �����]     ��       �� ���       ����
 � �����  �  u         ����  : ;           � ��       �����^  �   ��  	     �� ���       ����
 �����  �  u         ����  & '           +[ +]       ����.T  ��   	         �� ���        ����
 � �����  �  v         ����  ( )           1_ 1a       ����ZU  ު           �� ���        ����
 � �����  �  v         ����  * +           7c 7e       �����V  ·           �� ���        ����
 � �����  �  v         ����  , -           =g =i       �����W  ��           �� ���       ����
 � �����  �  v         ����  . /           Ck Cm       �����X  ��           �� ���       ����
 � �����  �  v         ����  0 1           Io Iq       ����
Z  n�           �� ���       ����
 � �����  �  v         ����  3 4           Os Ou       ����6[  R�           �� ���       ����
 � �����  �  v         ����  5 6           Uw Uy       ����b\  6�   ��       �� ���       ����
 � �����  �  v         ����  7 8           [{ [}       �����]     ��       �� ���       ����
 � �����  �  v         ����  9 :           a a�       �����^  �   ��  	     �� ���       ����
 �����  �  v         ����              � � [y       ����.T  ��   	   !      �� ���        ����
 � �����  �  w         ����               � � b}       ����ZU  ު      !     �� ���        ����
 � �����  �  w         ����  ! "           � � i�       �����V  ·      !     �� ���        ����
 � �����  �  w         ����  # $           � � p�       �����W  ��      !     �� ���       ����
 � �����  �  w         ����  % &           � � w�       �����X  ��      !     �� ���       ����
 � �����  �  w         ����  ' (           � � ~�       ����
Z  n�      !     �� ���       ����
 � �����  �  w         ����  ) *           � � ��       ����6[  R�      !     �� ���       ����
 � �����  �  w         ����  + ,           � � ��       ����b\  6�   ��  !     �� ���       ����
 � �����  �  w         ����  - .           � � ��       �����]     ��  !     �� ���       ����
 � �����  �  w         ����  / 0           � � ��       �����^  �   ��  !	     �� ���       ����
 �����  �  w         ����  3 4           r� h \       �����U  *�   	   N      �� ���        ����
 � �����  �  x         ����  5 6           y� l `       �����V  �      N     �� ���        ����
 � �����  �  x         ����  7 8           �� p d       ����X  ��      N     �� ���        ����
 � �����  �  x         ����  : ;           �� t h       ����BY  ��      N     �� ���       ����
 � �����  �  x         ����  < =           �� x l       ����nZ  ��      N     �� ���       ����
 � �����  �  x         ����  > ?           �� | p       �����[  ��      N     �� ���       ����
 � �����  �  x         ����  @ A           �� � t       �����\  ��      N     �� ���       ����
 � �����  �  x         ����  B C           �� � x       �����]  f	   ��  N     �� ���       ����
 � �����  �  x         ����  E F           �� � |       ����_  J   ��  N     �� ���       ����
 � �����  �  x         ����  G H           �� � �       ����J`  .#   ��  N	     �� ���       ����
 �����  �  x         ����  ' (           � � kb       �����U  *�   	   ]      �� ���        ����
 � �����  �  y         ����  ) *           � � rf       �����V  �      ]     �� ���        ����
 � �����  �  y         ����  + ,           � � yj       ����X  ��      ]     �� ���        ����
 � �����  �  y         ����  - .           � � �n       ����BY  ��      ]     �� ���       ����
 � �����  �  y         ����  / 0           � � �r       ����nZ  ��      ]     �� ���       ����
 � �����  �  y         ����  1 2           � � �v       �����[  ��      ]     �� ���       ����
 � �����  �  y         ����  4 5           � � �z       �����\  ��      ]     �� ���       ����
 � �����  �  y         ����  6 7           � � �~       �����]  f	   ��  ]     �� ���       ����
 � �����  �  y         ����  8 9           � ��       ����_  J   ��  ]     �� ���       ����
 � �����  �  y         ����  : ;           � ��       ����J`  .#   ��  ]	     �� ���       ����
 �����  �  y         ����  & '           .[ .]       �����U  *�   	   l      �� ���        ����
 � �����  �  z         ����  ( )           4_ 4a       �����V  �      l     �� ���        ����
 � �����  �  z         ����  * +           :c :e       ����X  ��      l     �� ���        ����
 � �����  �  z         ����  , -           @g @i       ����BY  ��      l     �� ���       ����
 � �����  �  z         ����  . /           Fk Fm       ����nZ  ��      l     �� ���       ����
 � �����  �  z         ����  0 1           Lo Lq       �����[  ��      l     �� ���       ����
 � �����  �  z         ����  3 4           Rs Ru       �����\  ��      l     �� ���       ����
 � �����  �  z         ����  5 6           Xw Xy       �����]  f	   ��  l     �� ���       ����
 � �����  �  z         ����  7 8           ^{ ^}       ����_  J   ��  l     �� ���       ����
 � �����  �  z         ����  9 :           d d�       ����J`  .#   ��  l	     �� ���       ����
 �����  �  z         ����              � � ^~       �����U  *�   	   {      �� ���        ����
 � �����  �  {         ����               � � e�       �����V  �      {     �� ���        ����
 � �����  �  {         ����  ! "           � � l�       ����X  ��      {     �� ���        ����
 � �����  �  {         ����  # $           � � s�       ����BY  ��      {     �� ���       ����
 � �����  �  {         ����  % &           � � z�       ����nZ  ��      {     �� ���       ����
 � �����  �  {         ����  ' (           � � ��       �����[  ��      {     �� ���       ����
 � �����  �  {         ����  ) *           � � ��       �����\  ��      {     �� ���       ����
 � �����  �  {         ����  + ,           � � ��       �����]  f	   ��  {     �� ���       ����
 � �����  �  {         ����  - .           � � ��       ����_  J   ��  {     �� ���       ����
 � �����  �  {         ����  / 0           � � ��       ����J`  .#   ��  {	     �� ���       ����
 �����  �  {          ��n ��                           �����  �        3      ��X ���        ������  ����������������        ��d ��  d                        �   �  �        /     ��T ���        ������  ����������������        ��e ��  d                        �   �  �        0     ��U ���        ������  ����������������        ��o ��d d                        �   �  �        1     ��V ���        ������  ����������������        ��p ��  3                        �����  �        2      ��W ���        ������  ����������������          �� � �2    ( ( ( (          >  �	        m       i   �    �������c   ������������|            �� � �2    ( ( ( (          z  n
        m      i   �    �������c   ������������|            �� � �2    ( ( ( (          �  "        m      i   �    �������c   ������������|            �� � �2    ( ( ( (          �  �        m      i   �   �������c   ������������|            �� � �2    ( ( ( (           .  �        m      i   �   �������c   ������������|            �� � �2    ( ( ( (       !   j  >        m      i   �   �������c   ������������|            �� � �2    ( ( ( (       #   �  �        m      i   �   �������c   ������������|            �� � �2    ( ( ( (       %   �  �        m      i   �   �������c   ������������|            �� � �2    ( ( ( (       '     Z        m      i   �   �������c   ������������|            �� � �2    ( ( ( (       )   Z          m 	     i   �   �������c   ������������|         ����    <          d d d d       #   �  �        &        ���        ����c   ������������}         ����   " ?          i i i i       %   �  �        &       ���        ����c   ������������}         ����   % B          n n n n       '     Z        &       ���        ����c   ������������}         ����   ( E          s s s s       )   Z          &       ���       ����c   ������������}         ����   + H          x x x x       *   �  �        &       ���       ����c   ������������}         ����   . K          } } } }       ,   �  v        &       ���       ����c   ������������}         ����   1 N          � � � �       .     *        &       ���       ����c   ������������}         ����   4 Q          � � � �       0   J  �        &       ���       ����c   ������������}         ����   7 T          � � � �       2   �  �        &       ���       ����c   ������������}         ����   : W          � � � �       3   �  F        &	       ���       ����c   ������������}         ����    <          d d d d       #   �  �        :        ���        ����c   ������������~         ����   " ?          i i i i       %   �  �        :       ���        ����c   ������������~         ����   % B          n n n n       '     Z        :       ���        ����c   ������������~         ����   ( E          s s s s       )   Z          :       ���       ����c   ������������~         ����   + H          x x x x       *   �  �        :       ���       ����c   ������������~         ����   . K          } } } }       ,   �  v        :       ���       ����c   ������������~         ����   1 N          � � � �       .     *        :       ���       ����c   ������������~         ����   4 Q          � � � �       0   J  �        :       ���       ����c   ������������~         ����   7 T          � � � �       2   �  �        :       ���       ����c   ������������~         ����   : W          � � � �       3   �  F        :	       ���       ����c   ������������~         ����    <          d d d d       #   �  �        N        ���        ����c   ������������         ����   " ?          i i i i       %   �  �        N       ���        ����c   ������������         ����   % B          n n n n       '     Z        N       ���        ����c   ������������         ����   ( E          s s s s       )   Z          N       ���       ����c   ������������         ����   + H          x x x x       *   �  �        N       ���       ����c   ������������         ����   . K          } } } }       ,   �  v        N       ���       ����c   ������������         ����   1 N          � � � �       .     *        N       ���       ����c   ������������         ����   4 Q          � � � �       0   J  �        N       ���       ����c   ������������         ����   7 T          � � � �       2   �  �        N       ���       ����c   ������������         ����   : W          � � � �       3   �  F        N	       ���       ����c   ������������         ����    <          d d d d       #   �  �        b        ���        ����c   �������������         ����   " ?          i i i i       %   �  �        b       ���        ����c   �������������         ����   % B          n n n n       '     Z        b       ���        ����c   �������������         ����   ( E          s s s s       )   Z          b       ���       ����c   �������������         ����   + H          x x x x       *   �  �        b       ���       ����c   �������������         ����   . K          } } } }       ,   �  v        b       ���       ����c   �������������         ����   1 N          � � � �       .     *        b       ���       ����c   �������������         ����   4 Q          � � � �       0   J  �        b       ���       ����c   �������������         ����   7 T          � � � �       2   �  �        b       ���       ����c   �������������         ����   : W          � � � �       3   �  F        b	       ���       ����c   �������������         ����� ��                            �����  �        ?      ��Y ���        ������  ����������������       ����� ��                          ����,  �  X           ��Z ���        ������  ����������������       ����� ��                          ����,  �  X           ��Z ���        ������  ����������������       ����� ��                          ����,  �  X           ��Z ���        ������  ����������������       ����� ��                          ����,  �  X            ��Z ���        ������  ����������������       ����� ��                          ����,  �  X     !      ��Z ���        ������  ����������������       ����� ��                          ����,  �  X     "      ��Z ���        ������  ����������������       ����� ��                       ;   ����,  �  X     #      ��[ ���        ������  ����������������       ����� ��                       ;   ����,  �  X     $      ��[ ���        ������  ����������������       ����� ��                       ;   ����,  �  X     %      ��[ ���        ������  ����������������       ����� ��                       ;   ����,  �  X     &      ��[ ���        ������  ����������������       ����� ��                       ;   ����,  �  X     '      ��[ ���        ������  ����������������       ����� ��                       ;   ����,  �  X     (      ��[ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     )      ��\ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     *      ��\ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     +      ��\ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     ,      ��\ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     -      ��\ ���        ������  ����������������       ����� ��                      < �   ����,  �  X     .      ��\ ���        ������  ����������������        ��s ��     
                    �����  �  [     4      ��] ���        ������  ����������������       ����� ��                            �����  �        @      ��^ ���        ������  ����������������        ��p ��  9                        �����  �        5      ��_ ���        ������  ����������������        ��p ��                           �����  �        6      ��` ���        ������  ����������������        ��o ��d d                        �����  �        7      ��a ���        ������  ����������������          �� � �2                    z  n
                   �    �������c   �������������            �� � �2      �              �  "                  �    �������c   �������������            �� � �2      �              �  �                  �    �������c   �������������            �� � �2      �               .  �                  �   �������c   �������������            �� � �2      �           !   j  >                  �   �������c   �������������            �� � �2      �           #   �  �                  �   �������c   �������������            �� � �2      �           %   �  �                  �   �������c   �������������            �� � �2      �           '     Z                  �   �������c   �������������            �� � �2      �           )   Z                    �   �������c   �������������            �� � �2      �           *   �  �         	         �   �������c   �������������            �� � �2        �         @   J  (        n       j   �    �������c   �������������            �� � �2        �         D   �  �        n      j   �    �������c   �������������            �� � �2        �         G   �  �        n      j   �    �������c   �������������            �� � �2        �         K   X  `        n      j   �   �������c   �������������            �� � �2        �         N   �  �        n      j   �   �������c   �������������            �� � �2        �         R     0         n      j   �   �������c   �������������            �� � �2        �         V   f  �!        n      j   �   �������c   �������������            �� � �2        �         Y   �   #        n      j   �   �������c   �������������            �� � �2        �         ]   	  h$        n      j   �   �������c   �������������            �� � �2        �         `   t	  �%        n 	     j   �   �������c   �������������              � �
2      J \            �  �        �       �   �    �������c   �������������              � �
2      L `             .  �        �      �   �    �������c   �������������              � �
2      N d         !   j  >        �      �   �    �������c   �������������              � �
2      P h         #   �  �        �      �   �   �������c   �������������              � �
2      R l         %   �  �        �      �   �   �������c   �������������              � �
2      T p         '     Z        �      �   �   �������c   �������������              � �
2      V t         )   Z          �      �   �   �������c   �������������              � �
2      X x         *   �  �        �      �   �   �������c   �������������              � �
2      Z |         ,   �  v        �      �   �   �������c   �������������              � �
2      \ �         .     *        � 	     �   �   �������c   �������������         ����    <          ( ( ( (       N   �  �        '        ���        ����c   �������������         ����    <          ( ( ( (       R     0         '       ���        ����c   �������������         ����    <          ( ( ( (       V   f  �!        '       ���        ����c   �������������         ����    <          ( ( ( (       Y   �   #        '       ���       ����c   �������������         ����    <          ( ( ( (       ]   	  h$        '       ���       ����c   �������������         ����    <          ( ( ( (       `   t	  �%        '       ���       ����c   �������������         ����    <          ( ( ( (       d   �	  8'        '       ���       ����c   �������������         ����    <          ( ( ( (       h   (
  �(        '       ���       ����c   �������������         ����    <          ( ( ( (       k   �
  *        '       ���       ����c   �������������         ����    <          ( ( ( (       o   �
  p+        '	       ���       ����c   �������������         ����    <          ( ( ( (       �   D  T=        (        ���        ����c   �������������         ����    <          ( ( ( (       �   �  �?        (       ���        ����c   �������������         ����    <          ( ( ( (       �   4  B        (       ���        ����c   �������������         ����    <          ( ( ( (       �   �  \D        (       ���       ����c   �������������         ����    <          ( ( ( (       �   $  �F        (       ���       ����c   �������������         ����    <          ( ( ( (       �   �  I        (       ���       ����c   �������������         ����    <          ( ( ( (       �     dK        (       ���       ����c   �������������         ����    <          ( ( ( (       �   �  �M        (       ���       ����c   �������������         ����    <          ( ( ( (       �     P        (       ���       ����c   �������������         ����    <          ( ( ( (       �   |  lR        (	       ���       ����c   �������������         ����    <          ( ( ( (       N   �  �        ;        ���        ����c   �������������         ����    <          ( ( ( (       R     0         ;       ���        ����c   �������������         ����    <          ( ( ( (       V   f  �!        ;       ���        ����c   �������������         ����    <          ( ( ( (       Y   �   #        ;       ���       ����c   �������������         ����    <          ( ( ( (       ]   	  h$        ;       ���       ����c   �������������         ����    <          ( ( ( (       `   t	  �%        ;       ���       ����c   �������������         ����    <          ( ( ( (       d   �	  8'        ;       ���       ����c   �������������         ����    <          ( ( ( (       h   (
  �(        ;       ���       ����c   �������������         ����    <          ( ( ( (       k   �
  *        ;       ���       ����c   �������������         ����    <          ( ( ( (       o   �
  p+        ;	       ���       ����c   �������������         ����    <          ( ( ( (       �   D  T=        <        ���        ����c   �������������         ����    <          ( ( ( (       �   �  �?        <       ���        ����c   �������������         ����    <          ( ( ( (       �   4  B        <       ���        ����c   �������������         ����    <          ( ( ( (       �   �  \D        <       ���       ����c   �������������         ����    <          ( ( ( (       �   $  �F        <       ���       ����c   �������������         ����    <          ( ( ( (       �   �  I        <       ���       ����c   �������������         ����    <          ( ( ( (       �     dK        <       ���       ����c   �������������         ����    <          ( ( ( (       �   �  �M        <       ���       ����c   �������������         ����    <          ( ( ( (       �     P        <       ���       ����c   �������������         ����    <          ( ( ( (       �   |  lR        <	       ���       ����c   �������������         ����    <          ( ( ( (       N   �  �        O        ���        ����c   �������������         ����    <          ( ( ( (       R     0         O       ���        ����c   �������������         ����    <          ( ( ( (       V   f  �!        O       ���        ����c   �������������         ����    <          ( ( ( (       Y   �   #        O       ���       ����c   �������������         ����    <          ( ( ( (       ]   	  h$        O       ���       ����c   �������������         ����    <          ( ( ( (       `   t	  �%        O       ���       ����c   �������������         ����    <          ( ( ( (       d   �	  8'        O       ���       ����c   �������������         ����    <          ( ( ( (       h   (
  �(        O       ���       ����c   �������������         ����    <          ( ( ( (       k   �
  *        O       ���       ����c   �������������         ����    <          ( ( ( (       o   �
  p+        O	       ���       ����c   �������������         ����    <          ( ( ( (       �   D  T=        P        ���        ����c   �������������         ����    <          ( ( ( (       �   �  �?        P       ���        ����c   �������������         ����    <          ( ( ( (       �   4  B        P       ���        ����c   �������������         ����    <          ( ( ( (       �   �  \D        P       ���       ����c   �������������         ����    <          ( ( ( (       �   $  �F        P       ���       ����c   �������������         ����    <          ( ( ( (       �   �  I        P       ���       ����c   �������������         ����    <          ( ( ( (       �     dK        P       ���       ����c   �������������         ����    <          ( ( ( (       �   �  �M        P       ���       ����c   �������������         ����    <          ( ( ( (       �     P        P       ���       ����c   �������������         ����    <          ( ( ( (       �   |  lR        P	       ���       ����c   �������������         ����    <          ( ( ( (       N   �  �        c        ���        ����c   �������������         ����    <          ( ( ( (       R     0         c       ���        ����c   �������������         ����    <          ( ( ( (       V   f  �!        c       ���        ����c   �������������         ����    <          ( ( ( (       Y   �   #        c       ���       ����c   �������������         ����    <          ( ( ( (       ]   	  h$        c       ���       ����c   �������������         ����    <          ( ( ( (       `   t	  �%        c       ���       ����c   �������������         ����    <          ( ( ( (       d   �	  8'        c       ���       ����c   �������������         ����    <          ( ( ( (       h   (
  �(        c       ���       ����c   �������������         ����    <          ( ( ( (       k   �
  *        c       ���       ����c   �������������         ����    <          ( ( ( (       o   �
  p+        c	       ���       ����c   �������������         ����    <          ( ( ( (       �   D  T=        d        ���        ����c   �������������         ����    <          ( ( ( (       �   �  �?        d       ���        ����c   �������������         ����    <          ( ( ( (       �   4  B        d       ���        ����c   �������������         ����    <          ( ( ( (       �   �  \D        d       ���       ����c   �������������         ����    <          ( ( ( (       �   $  �F        d       ���       ����c   �������������         ����    <          ( ( ( (       �   �  I        d       ���       ����c   �������������         ����    <          ( ( ( (       �     dK        d       ���       ����c   �������������         ����    <          ( ( ( (       �   �  �M        d       ���       ����c   �������������         ����    <          ( ( ( (       �     P        d       ���       ����c   �������������         ����    <          ( ( ( (       �   |  lR        d	       ���       ����c   �������������         ����  2 3          _� h \       �  �M  :Y   	   �      �   �        ����
 � �����  �  �         ����  4 5          f� l `       �  O  f      �     �   �        ����
 � �����  �  �         ����  6 7          m� p d       �  FP  s      �     �   �        ����
 � �����  �  �         ����  9 :          t� t h       �  rQ  �      �     �   �       ����
 � �����  �  �         ����  ; <          {� x l       	  �R  ʌ      �     �   �       ����
 � �����  �  �         ����  = >          �� | p       7	  �S  ��      �     �   �       ����
 � �����  �  �         ����  ? @          �� � t       X	  �T  ��      �     �   �       ����
 � �����  �  �         ����  A B          �� � x       y	  "V  v�   ��  �     �   �       ����
 � �����  �  �         ����  D E          �� � |       �	  NW  Z�   ��  �     �   �       ����
 � �����  �  �         ����  F G          �� � �       �	  zX  >�   ��  �	     �   �       ����
 7  �  �  �         ����  ' (          � � Xb       �  �M  :Y   	   �      �   �        ����
 � �����  �  �         ����  ) *          � � _f       �  O  f      �     �   �        ����
 � �����  �  �         ����  + ,          � � fj       �  FP  s      �     �   �        ����
 � �����  �  �         ����  - .          � � mn       �  rQ  �      �     �   �       ����
 � �����  �  �         ����  / 0          � � tr       	  �R  ʌ      �     �   �       ����
 � �����  �  �         ����  1 2          � � {v       7	  �S  ��      �     �   �       ����
 � �����  �  �         ����  4 5          � � �z       X	  �T  ��      �     �   �       ����
 � �����  �  �         ����  6 7          � � �~       y	  "V  v�   ��  �     �   �       ����
 � �����  �  �         ����  8 9          � � ��       �	  NW  Z�   ��  �     �   �       ����
 � �����  �  �         ����  : ;          � � ��       �	  zX  >�   ��  �	     �   �       ����
 7  �  �  �         ����  & '          [ ]       �  �M  :Y   	   �      �   �        ����
 � �����  �  �         ����  ( )          !_ !a       �  O  f      �     �   �        ����
 � �����  �  �         ����  * +          'c 'e       �  FP  s      �     �   �        ����
 � �����  �  �         ����  , -          -g -i       �  rQ  �      �     �   �       ����
 � �����  �  �         ����  . /          3k 3m       	  �R  ʌ      �     �   �       ����
 � �����  �  �         ����  0 1          9o 9q       7	  �S  ��      �     �   �       ����
 � �����  �  �         ����  3 4          ?s ?u       X	  �T  ��      �     �   �       ����
 � �����  �  �         ����  5 6          Ew Ey       y	  "V  v�   ��  �     �   �       ����
 � �����  �  �         ����  7 8          K{ K}       �	  NW  Z�   ��  �     �   �       ����
 � �����  �  �         ����  9 :          Q Q�       �	  zX  >�   ��  �	     �   �       ����
 7  �  �  �         ����   7 8          �� v j d     n
  �V  �               ���        ���� � �����  �  �         ����   9 :          �� { o e     �
  4X  p"              ���        ���� � �����  �  �         ����   ; <          �� � t f     �
  ~Y  �1              ���        ���� � �����  �  �         ����   > ?          �� � y g     �
  �Z  `A              ���       ���� � �����  �  �         ����   @ A          �� � ~ h       \  �P              ���       ���� � �����  �  �         ����   B C          �� � � i     4  \]  P`   ��          ���       ���� � �����  �  �         ����   D E          �� � j     [  �^  �o   ��          ���       ���� � �����  �  �         ����   F G          �� � k     �  �_  @   ��          ���       ���� � �����  �  �         ����   I J          �� � l     �  :a  ��   ��          ���       ���� �����  �  �         ����   K L          �� � m     �  �b  0�   ��   	       ���       ���� A  �  �  �         ����   + ,          � � zp d     n
  �V  �      4        ���        ���� � �����  �  �         ����   - .          � � �u e     �
  4X  p"      4       ���        ���� � �����  �  �         ����   / 0          � � �z f     �
  ~Y  �1      4       ���        ���� � �����  �  �         ����   1 2          � � � g     �
  �Z  `A      4       ���       ���� � �����  �  �         ����   3 4          � � �� h       \  �P      4       ���       ���� � �����  �  �         ����   5 6          � � �� i     4  \]  P`   ��  4       ���       ���� � �����  �  �         ����   8 9          � � �� j     [  �^  �o   ��  4       ���       ���� � �����  �  �         ����   : ;          � �� k     �  �_  @   ��  4       ���       ���� � �����  �  �         ����   < =          � �� l     �  :a  ��   ��  4       ���       ���� �����  �  �         ����   > ?          � �� m     �  �b  0�   ��  4	       ���       ���� A  �  �  �         ����   * +          5i 5k d     n
  �V  �      H        ���        ���� � �����  �  �         ����   , -          <n <p e     �
  4X  p"      H       ���        ���� � �����  �  �         ����   . /          Cs Cu f     �
  ~Y  �1      H       ���        ���� � �����  �  �         ����   0 1          Jx Jz g     �
  �Z  `A      H       ���       ���� � �����  �  �         ����   2 3          Q} Q h       \  �P      H       ���       ���� � �����  �  �         ����   4 5          X� X� i     4  \]  P`   ��  H       ���       ���� � �����  �  �         ����   7 8          _� _� j     [  �^  �o   ��  H       ���       ���� � �����  �  �         ����   9 :          f� f� k     �  �_  @   ��  H       ���       ���� � �����  �  �         ����   ; <          m� m� l     �  :a  ��   ��  H       ���       ���� �����  �  �         ����   = >          t� t� m     �  �b  0�   ��  H	       ���       ���� A  �  �  �         ����     !          � � |q d     n
  �V  �      \        ���        ���� � �����  �  �         ����   " #          � � �v e     �
  4X  p"      \       ���        ���� � �����  �  �         ����   $ %          � � �{ f     �
  ~Y  �1      \       ���        ���� � �����  �  �         ����   & '          � � �� g     �
  �Z  `A      \       ���       ���� � �����  �  �         ����   ( )          � � �� h       \  �P      \       ���       ���� � �����  �  �         ����   * +          � � �� i     4  \]  P`   ��  \       ���       ���� � �����  �  �         ����   , -          � � �� j     [  �^  �o   ��  \       ���       ���� � �����  �  �         ����   . /          � � �� k     �  �_  @   ��  \       ���       ���� � �����  �  �         ����   0 1          � � �� l     �  :a  ��   ��  \       ���       ���� �����  �  �         ����   2 3          � �� m     �  �b  0�   ��  \	       ���       ���� A  �  �  �         ����  5 6          l� v j d     2
  �T  ��      �        ���        ���� � �����  �  �         ����  7 8          s� { o e     Y
  @V         �       ���        ���� � �����  �  �         ����  9 :          z� � t f     �
  �W  x      �       ���        ���� � �����  �  �         ����  < =          �� � y g     �
  �X  �)      �       ���       ���� � �����  �  �         ����  > ?          �� � ~ h     �
  Z  h9      �       ���       ���� � �����  �  �         ����  @ A          �� � � i     �
  h[  �H   ��  �       ���       ���� � �����  �  �         ����  B C          �� � j       �\  XX   ��  �       ���       ���� � �����  �  �         ����  D E          �� � k     G  �]  �g   ��  �       ���       ���� � �����  �  �         ����  G H          �� � l     n  F_  Hw   ��  �       ���       ���� �����  �  �         ����  I J          �� � m     �  �`  ��   ��  �	       ���       ���� A  �  �  �         ����  * +          � � ep d     2
  �T  ��      �        ���        ���� � �����  �  �         ����  , -          � � lu e     Y
  @V         �       ���        ���� � �����  �  �         ����  . /          � � sz f     �
  �W  x      �       ���        ���� � �����  �  �         ����  0 1          � � z g     �
  �X  �)      �       ���       ���� � �����  �  �         ����  2 3          � � �� h     �
  Z  h9      �       ���       ���� � �����  �  �         ����  4 5          � � �� i     �
  h[  �H   ��  �       ���       ���� � �����  �  �         ����  7 8          � � �� j       �\  XX   ��  �       ���       ���� � �����  �  �         ����  9 :          � � �� k     G  �]  �g   ��  �       ���       ���� � �����  �  �         ����  ; <          � � �� l     n  F_  Hw   ��  �       ���       ���� �����  �  �         ����  = >          � � �� m     �  �`  ��   ��  �	       ���       ���� A  �  �  �         ����  ) *           i  k d     2
  �T  ��      �        ���        ���� � �����  �  �         ����  + ,          'n 'p e     Y
  @V         �       ���        ���� � �����  �  �         ����  - .          .s .u f     �
  �W  x      �       ���        ���� � �����  �  �         ����  / 0          5x 5z g     �
  �X  �)      �       ���       ���� � �����  �  �         ����  1 2          <} < h     �
  Z  h9      �       ���       ���� � �����  �  �         ����  3 4          C� C� i     �
  h[  �H   ��  �       ���       ���� � �����  �  �         ����  6 7          J� J� j       �\  XX   ��  �       ���       ���� � �����  �  �         ����  8 9          Q� Q� k     G  �]  �g   ��  �       ���       ���� � �����  �  �         ����  : ;          X� X� l     n  F_  Hw   ��  �       ���       ���� �����  �  �         ����  < =          _� _� m     �  �`  ��   ��  �	       ���       ���� A  �  �  �         ����              � � sh d     2
  �T  ��      �        ���        ���� � �����  �  �         ����  ! "          � � zm e     Y
  @V         �       ���        ���� � �����  �  �         ����  # $          � � �r f     �
  �W  x      �       ���        ���� � �����  �  �         ����  % &          � � �w g     �
  �X  �)      �       ���       ���� � �����  �  �         ����  ' (          � � �| h     �
  Z  h9      �       ���       ���� � �����  �  �         ����  ) *          � � �� i     �
  h[  �H   ��  �       ���       ���� � �����  �  �         ����  + ,          � � �� j       �\  XX   ��  �       ���       ���� � �����  �  �         ����  - .          � � �� k     G  �]  �g   ��  �       ���       ���� � �����  �  �         ����  / 0          � � �� l     n  F_  Hw   ��  �       ���       ���� �����  �  �         ����  1 2          � � �� m     �  �`  ��   ��  �	       ���       ���� A  �  �  �          ��  8 9           �� v j �     �����^  �p       �       �    �        ���� � �����  �  �          ��  : ;           �� { o �     ����`  0�       �      �    �        ���� � �����  �  �          ��  < =           �� � t �     ����Na  ��       �      �    �        ���� � �����  �  �          ��  ? @           �� � y �     �����b   �       �      �    �        ���� � �����  �  �          ��  A B           �� � ~ �     �����c  ��       �      �    �        ���� � �����  �  �          ��  C D           �� � � �     ����,e  �       �      �    �        ���� � �����  �  �          ��  E F           �� � �     ����vf  ��       �      �    �        ���� � �����  �  �          ��  G H           �� � �     �����g   �       �      �    �        ���� � �����  �  �          ��  J K           �� � �     ����
i  x�       �      �    �        ���� �����  �  �          ��  L M           �� � �     ����Tj  ��       � 	     �    �        ���� �����  �  �          ��  + ,           � � �p �     �����^  �p       �       �    �        ���� � �����  �  �          ��  - .           � � �u �     ����`  0�       �      �    �        ���� � �����  �  �          ��  / 0           � � �z �     ����Na  ��       �      �    �        ���� � �����  �  �          ��  1 2           � � � �     �����b   �       �      �    �        ���� � �����  �  �          ��  3 4           � �� �     �����c  ��       �      �    �        ���� � �����  �  �          ��  5 6           � �� �     ����,e  �       �      �    �        ���� � �����  �  �          ��  8 9           � �� �     ����vf  ��       �      �    �        ���� � �����  �  �          ��  : ;           � �� �     �����g   �       �      �    �        ���� � �����  �  �          ��  < =           � �� �     ����
i  x�       �      �    �        ���� �����  �  �          ��  > ?           �  �� �     ����Tj  ��       � 	     �    �        ���� �����  �  �          ��  * +           Gi Gk �     �����^  �p       �       �    �        ���� � �����  �  �          ��  , -           Nn Np �     ����`  0�       �      �    �        ���� � �����  �  �          ��  . /           Us Uu �     ����Na  ��       �      �    �        ���� � �����  �  �          ��  0 1           \x \z �     �����b   �       �      �    �        ���� � �����  �  �          ��  2 3           c} c �     �����c  ��       �      �    �        ���� � �����  �  �          ��  4 5           j� j� �     ����,e  �       �      �    �        ���� � �����  �  �          ��  7 8           q� q� �     ����vf  ��       �      �    �        ���� � �����  �  �          ��  9 :           x� x� �     �����g   �       �      �    �        ���� � �����  �  �          ��  ; <           � � �     ����
i  x�       �      �    �        ���� �����  �  �          ��  = >           �� �� �     ����Tj  ��       � 	     �    �        ���� �����  �  �          ��    !           � � � �     �����^  �p       �       �    �        ���� � �����  �  �          ��  " #           � � �� �     ����`  0�       �      �    �        ���� � �����  �  �          ��  $ %           � � �� �     ����Na  ��       �      �    �        ���� � �����  �  �          ��  & '           � � �� �     �����b   �       �      �    �        ���� � �����  �  �          ��  ( )           � � �� �     �����c  ��       �      �    �        ���� � �����  �  �          ��  * +           � � �� �     ����,e  �       �      �    �        ���� � �����  �  �          ��  , -           � � �� �     ����vf  ��       �      �    �        ���� � �����  �  �          ��  . /           � � �� �     �����g   �       �      �    �        ���� � �����  �  �          ��  0 1           � �� �     ����
i  x�       �      �    �        ���� �����  �  �          ��  2 3           � �� �     ����Tj  ��       � 	     �    �        ���� �����  �  �         ����  6 7          y� v j d     &
  �T  ��      �        ���        ���� � �����  �  �         ����  8 9          �� { o e     M
  �U  P      �       ���        ���� � �����  �  �         ����  : ;          �� � t f     u
  &W  �      �       ���        ���� � �����  �  �         ����  = >          �� � y g     �
  pX  @%      �       ���       ���� � �����  �  �         ����  ? @          �� � ~ h     �
  �Y  �4      �       ���       ���� � �����  �  �         ����  A B          �� � � i     �
  [  0D   ��  �       ���       ���� � �����  �  �         ����  C D          �� � j       N\  �S   ��  �       ���       ���� � �����  �  �         ����  E F          �� � k     ;  �]   c   ��  �       ���       ���� � �����  �  �         ����  H I          �� � l     b  �^  �r   ��  �       ���       ���� �����  �  �         ����  J K          �� � m     �  ,`  �   ��  �	       ���       ���� A  �  �  �         ����  * +          � � rp d     &
  �T  ��              ���        ���� � �����  �  �         ����  , -          � � yu e     M
  �U  P             ���        ���� � �����  �  �         ����  . /          � � �z f     u
  &W  �             ���        ���� � �����  �  �         ����  0 1          � � � g     �
  pX  @%             ���       ���� � �����  �  �         ����  2 3          � � �� h     �
  �Y  �4             ���       ���� � �����  �  �         ����  4 5          � � �� i     �
  [  0D   ��         ���       ���� � �����  �  �         ����  7 8          � � �� j       N\  �S   ��         ���       ���� � �����  �  �         ����  9 :          � � �� k     ;  �]   c   ��         ���       ���� � �����  �  �         ����  ; <          �  �� l     b  �^  �r   ��         ���       ���� �����  �  �         ����  = >          � �� m     �  ,`  �   ��  	       ���       ���� A  �  �  �         ����  ) *          -i -k d     &
  �T  ��              ���        ���� � �����  �  �         ����  + ,          4n 4p e     M
  �U  P             ���        ���� � �����  �  �         ����  - .          ;s ;u f     u
  &W  �             ���        ���� � �����  �  �         ����  / 0          Bx Bz g     �
  pX  @%             ���       ���� � �����  �  �         ����  1 2          I} I h     �
  �Y  �4             ���       ���� � �����  �  �         ����  3 4          P� P� i     �
  [  0D   ��         ���       ���� � �����  �  �         ����  6 7          W� W� j       N\  �S   ��         ���       ���� � �����  �  �         ����  8 9          ^� ^� k     ;  �]   c   ��         ���       ���� � �����  �  �         ����  : ;          e� e� l     b  �^  �r   ��         ���       ���� �����  �  �         ����  < =          l� l� m     �  ,`  �   ��  	       ���       ���� A  �  �  �         ����              � � vq d     &
  �T  ��      -        ���        ���� � �����  �  �         ����  ! "          � � }v e     M
  �U  P      -       ���        ���� � �����  �  �         ����  # $          � � �{ f     u
  &W  �      -       ���        ���� � �����  �  �         ����  % &          � � �� g     �
  pX  @%      -       ���       ���� � �����  �  �         ����  ' (          � � �� h     �
  �Y  �4      -       ���       ���� � �����  �  �         ����  ) *          � � �� i     �
  [  0D   ��  -       ���       ���� � �����  �  �         ����  + ,          � � �� j       N\  �S   ��  -       ���       ���� � �����  �  �         ����  - .          � � �� k     ;  �]   c   ��  -       ���       ���� � �����  �  �         ����  / 0          � � �� l     b  �^  �r   ��  -       ���       ���� �����  �  �         ����  1 2          � �� m     �  ,`  �   ��  -	       ���       ���� A  �  �  �         ����  5 6          g� v j d     �
  �[  8K      `        ���        ���� � �����  �  �         ����  7 8          n� { o e     %  �\  �Z      `       ���        ���� � �����  �  �         ����  9 :          u� � t f     M  .^  (j      `       ���        ���� � �����  �  �         ����  < =          |� � y g     t  x_  �y      `       ���       ���� � �����  �  �         ����  > ?          �� � ~ h     �  �`  �      `       ���       ���� � �����  �  �         ����  @ A          �� � � i     �  b  ��   ��  `       ���       ���� � �����  �  �         ����  B C          �� � j     �  Vc  �   ��  `       ���       ���� � �����  �  �         ����  D E          �� � k       �d  ��   ��  `       ���       ���� � �����  �  �         ����  G H          �� � l     :  �e  ��   ��  `       ���       ���� �����  �  �         ����  I J          �� � m     b  4g  p�   ��  `	       ���       ���� A  �  �  �         ����  * +          � � `p d     �
  �[  8K      q        ���        ���� � �����  �  �         ����  , -          � � gu e     %  �\  �Z      q       ���        ���� � �����  �  �         ����  . /          � � nz f     M  .^  (j      q       ���        ���� � �����  �  �         ����  0 1          � � u g     t  x_  �y      q       ���       ���� � �����  �  �         ����  2 3          � � |� h     �  �`  �      q       ���       ���� � �����  �  �         ����  4 5          � � �� i     �  b  ��   ��  q       ���       ���� � �����  �  �         ����  7 8          � � �� j     �  Vc  �   ��  q       ���       ���� � �����  �  �         ����  9 :          � � �� k       �d  ��   ��  q       ���       ���� � �����  �  �         ����  ; <          � � �� l     :  �e  ��   ��  q       ���       ���� �����  �  �         ����  = >          � � �� m     b  4g  p�   ��  q	       ���       ���� A  �  �  �         ����  ) *          i k d     �
  �[  8K      �        ���        ���� � �����  �  �         ����  + ,          "n "p e     %  �\  �Z      �       ���        ���� � �����  �  �         ����  - .          )s )u f     M  .^  (j      �       ���        ���� � �����  �  �         ����  / 0          0x 0z g     t  x_  �y      �       ���       ���� � �����  �  �         ����  1 2          7} 7 h     �  �`  �      �       ���       ���� � �����  �  �         ����  3 4          >� >� i     �  b  ��   ��  �       ���       ���� � �����  �  �         ����  6 7          E� E� j     �  Vc  �   ��  �       ���       ���� � �����  �  �         ����  8 9          L� L� k       �d  ��   ��  �       ���       ���� � �����  �  �         ����  : ;          S� S� l     :  �e  ��   ��  �       ���       ���� �����  �  �         ����  < =          Z� Z� m     b  4g  p�   ��  �	       ���       ���� A  �  �  �         ����              } � pe d     �
  �[  8K      �        ���        ���� � �����  �  �         ����  ! "          � � wj e     %  �\  �Z      �       ���        ���� � �����  �  �         ����  # $          � � ~o f     M  .^  (j      �       ���        ���� � �����  �  �         ����  % &          � � �t g     t  x_  �y      �       ���       ���� � �����  �  �         ����  ' (          � � �y h     �  �`  �      �       ���       ���� � �����  �  �         ����  ) *          � � �~ i     �  b  ��   ��  �       ���       ���� � �����  �  �         ����  + ,          � � �� j     �  Vc  �   ��  �       ���       ���� � �����  �  �         ����  - .          � � �� k       �d  ��   ��  �       ���       ���� � �����  �  �         ����  / 0          � � �� l     :  �e  ��   ��  �       ���       ���� �����  �  �         ����  1 2          � � �� m     b  4g  p�   ��  �	       ���       ���� A  �  �  �         ����  8 9          �� v j d     �
  
Z  x8      �      
  ���        ���� � �����  �  �         ����  : ;          �� { o e     �
  T[  �G      �     
  ���        ���� � �����  �  �         ����  < =          �� � t f       �\  hW      �     
  ���        ���� � �����  �  �         ����  ? @          �� � y g     D  �]  �f      �     
  ���       ���� � �����  �  �         ����  A B          �� � ~ h     l  2_  Xv      �     
  ���       ���� � �����  �  �         ����  C D          �� � � i     �  |`  Ѕ   ��  �     
  ���       ���� � �����  �  �         ����  E F          �� � j     �  �a  H�   ��  �     
  ���       ���� � �����  �  �         ����  G H          �� � k     �  c  ��   ��  �     
  ���       ���� � �����  �  �         ����  J K          �� � l     
  Zd  8�   ��  �     
  ���       ���� �����  �  �         ����  L M          �� � m     2  �e  ��   ��  �	     
  ���       ���� A  �  �  �         ����  + ,          � � �p d     �
  
Z  x8      �      
  ���        ���� � �����  �  �         ����  - .          � � �u e     �
  T[  �G      �     
  ���        ���� � �����  �  �         ����  / 0          � � �z f       �\  hW      �     
  ���        ���� � �����  �  �         ����  1 2          � � � g     D  �]  �f      �     
  ���       ���� � �����  �  �         ����  3 4          � � �� h     l  2_  Xv      �     
  ���       ���� � �����  �  �         ����  5 6          � �� i     �  |`  Ѕ   ��  �     
  ���       ���� � �����  �  �         ����  8 9          � 	�� j     �  �a  H�   ��  �     
  ���       ���� � �����  �  �         ����  : ;          � �� k     �  c  ��   ��  �     
  ���       ���� � �����  �  �         ����  < =          � �� l     
  Zd  8�   ��  �     
  ���       ���� �����  �  �         ����  > ?          � �� m     2  �e  ��   ��  �	     
  ���       ���� A  �  �  �         ����  * +          Bi Bk d     �
  
Z  x8      �      
  ���        ���� � �����  �  �         ����  , -          In Ip e     �
  T[  �G      �     
  ���        ���� � �����  �  �         ����  . /          Ps Pu f       �\  hW      �     
  ���        ���� � �����  �  �         ����  0 1          Wx Wz g     D  �]  �f      �     
  ���       ���� � �����  �  �         ����  2 3          ^} ^ h     l  2_  Xv      �     
  ���       ���� � �����  �  �         ����  4 5          e� e� i     �  |`  Ѕ   ��  �     
  ���       ���� � �����  �  �         ����  7 8          l� l� j     �  �a  H�   ��  �     
  ���       ���� � �����  �  �         ����  9 :          s� s� k     �  c  ��   ��  �     
  ���       ���� � �����  �  �         ����  ; <          z� z� l     
  Zd  8�   ��  �     
  ���       ���� �����  �  �         ����  = >          �� �� m     2  �e  ��   ��  �	     
  ���       ���� A  �  �  �         ����    !          � � �� d     �
  
Z  x8      �      
  ���        ���� � �����  �  �         ����  " #          � � �� e     �
  T[  �G      �     
  ���        ���� � �����  �  �         ����  $ %          � � �� f       �\  hW      �     
  ���        ���� � �����  �  �         ����  & '          � � �� g     D  �]  �f      �     
  ���       ���� � �����  �  �         ����  ( )          � � �� h     l  2_  Xv      �     
  ���       ���� � �����  �  �         ����  * +          � � �� i     �  |`  Ѕ   ��  �     
  ���       ���� � �����  �  �         ����  , -          �  �� j     �  �a  H�   ��  �     
  ���       ���� � �����  �  �         ����  . /          � �� k     �  c  ��   ��  �     
  ���       ���� � �����  �  �         ����  0 1          � �� l     
  Zd  8�   ��  �     
  ���       ���� �����  �  �         ����  2 3          � �� m     2  �e  ��   ��  �	     
  ���       ���� A  �  �  �         ����  6 7          t� v j d     �
  zX  �%      ,        ���        ���� � �����  �  �         ����  8 9          {� { o e     �
  �Y  05      ,       ���        ���� � �����  �  �         ����  : ;          �� � t f     �
  [  �D      ,       ���        ���� � �����  �  �         ����  = >          �� � y g       X\   T      ,       ���       ���� � �����  �  �         ����  ? @          �� � ~ h     <  �]  �c      ,       ���       ���� � �����  �  �         ����  A B          �� � � i     d  �^  s   ��  ,       ���       ���� � �����  �  �         ����  C D          �� � j     �  6`  ��   ��  ,       ���       ���� � �����  �  �         ����  E F          �� � k     �  �a   �   ��  ,       ���       ���� � �����  �  �         ����  H I          �� � l     �  �b  x�   ��  ,       ���       ���� �����  �  �         ����  J K          �� � m       d  �   ��  ,	       ���       ���� A  �  �  �         ����  * +          � � mp d     �
  zX  �%      =        ���        ���� � �����  �  �         ����  , -          � � tu e     �
  �Y  05      =       ���        ���� � �����  �  �         ����  . /          � � {z f     �
  [  �D      =       ���        ���� � �����  �  �         ����  0 1          � � � g       X\   T      =       ���       ���� � �����  �  �         ����  2 3          � � �� h     <  �]  �c      =       ���       ���� � �����  �  �         ����  4 5          � � �� i     d  �^  s   ��  =       ���       ���� � �����  �  �         ����  7 8          � � �� j     �  6`  ��   ��  =       ���       ���� � �����  �  �         ����  9 :          � � �� k     �  �a   �   ��  =       ���       ���� � �����  �  �         ����  ; <          � � �� l     �  �b  x�   ��  =       ���       ���� �����  �  �         ����  = >          � �� m       d  �   ��  =	       ���       ���� A  �  �  �         ����  ) *          (i (k d     �
  zX  �%      N        ���        ���� � �����  �  �         ����  + ,          /n /p e     �
  �Y  05      N       ���        ���� � �����  �  �         ����  - .          6s 6u f     �
  [  �D      N       ���        ���� � �����  �  �         ����  / 0          =x =z g       X\   T      N       ���       ���� � �����  �  �         ����  1 2          D} D h     <  �]  �c      N       ���       ���� � �����  �  �         ����  3 4          K� K� i     d  �^  s   ��  N       ���       ���� � �����  �  �         ����  6 7          R� R� j     �  6`  ��   ��  N       ���       ���� � �����  �  �         ����  8 9          Y� Y� k     �  �a   �   ��  N       ���       ���� � �����  �  �         ����  : ;          `� `� l     �  �b  x�   ��  N       ���       ���� �����  �  �         ����  < =          g� g� m       d  �   ��  N	       ���       ���� A  �  �  �         ����              � � �w d     �
  zX  �%      _        ���        ���� � �����  �  �         ����  ! "          � � �| e     �
  �Y  05      _       ���        ���� � �����  �  �         ����  # $          � � �� f     �
  [  �D      _       ���        ���� � �����  �  �         ����  % &          � � �� g       X\   T      _       ���       ���� � �����  �  �         ����  ' (          � � �� h     <  �]  �c      _       ���       ���� � �����  �  �         ����  ) *          � � �� i     d  �^  s   ��  _       ���       ���� � �����  �  �         ����  + ,          � � �� j     �  6`  ��   ��  _       ���       ���� � �����  �  �         ����  - .          � � �� k     �  �a   �   ��  _       ���       ���� � �����  �  �         ����  / 0          � �� l     �  �b  x�   ��  _       ���       ���� �����  �  �         ����  1 2          � 	�� m       d  �   ��  _	       ���       ���� A  �  �  �         ����  7 8          �� v j d     .  *]  �]      �      �   �        ���� � �����  �  �         ����  9 :          �� { o e     U  t^  pm      �     �   �        ���� � �����  �  �         ����  ; <          �� � t f     }  �_  �|      �     �   �        ���� � �����  �  �         ����  > ?          �� � y g     �  a  `�      �     �   �       ���� � �����  �  �         ����  @ A          �� � ~ h     �  Rb  ؛      �     �   �       ���� � �����  �  �         ����  B C          �� � � i     �  �c  P�   ��  �     �   �       ���� � �����  �  �         ����  D E          �� � j       �d  Ⱥ   ��  �     �   �       ���� � �����  �  �         ����  F G          �� � k     C  0f  @�   ��  �     �   �       ���� � �����  �  �         ����  I J          �� � l     j  zg  ��   ��  �     �   �       ���� �����  �  �         ����  K L          �� � m     �  �h  0�   ��  �	     �   �       ���� A  �  �  �         ����  + ,          � � p d     .  *]  �]      �      �   �        ���� � �����  �  �         ����  - .          � � �u e     U  t^  pm      �     �   �        ���� � �����  �  �         ����  / 0          � � �z f     }  �_  �|      �     �   �        ���� � �����  �  �         ����  1 2          � � � g     �  a  `�      �     �   �       ���� � �����  �  �         ����  3 4          � � �� h     �  Rb  ؛      �     �   �       ���� � �����  �  �         ����  5 6          � � �� i     �  �c  P�   ��  �     �   �       ���� � �����  �  �         ����  8 9          � �� j       �d  Ⱥ   ��  �     �   �       ���� � �����  �  �         ����  : ;          � �� k     C  0f  @�   ��  �     �   �       ���� � �����  �  �         ����  < =          � �� l     j  zg  ��   ��  �     �   �       ���� �����  �  �         ����  > ?          � �� m     �  �h  0�   ��  �	     �   �       ���� A  �  �  �         ����  * +          :i :k d     .  *]  �]      �      �   �        ���� � �����  �  �         ����  , -          An Ap e     U  t^  pm      �     �   �        ���� � �����  �  �         ����  . /          Hs Hu f     }  �_  �|      �     �   �        ���� � �����  �  �         ����  0 1          Ox Oz g     �  a  `�      �     �   �       ���� � �����  �  �         ����  2 3          V} V h     �  Rb  ؛      �     �   �       ���� � �����  �  �         ����  4 5          ]� ]� i     �  �c  P�   ��  �     �   �       ���� � �����  �  �         ����  7 8          d� d� j       �d  Ⱥ   ��  �     �   �       ���� � �����  �  �         ����  9 :          k� k� k     C  0f  @�   ��  �     �   �       ���� � �����  �  �         ����  ; <          r� r� l     j  zg  ��   ��  �     �   �       ���� �����  �  �         ����  = >          y� y� m     �  �h  0�   ��  �	     �   �       ���� A  �  �  �         ����	  5 6           o� v j d     �����a  8�      �      �� ���        ���� � �����  �  �         ����	  7 8           v� { o e     ����$c  ��      �     �� ���        ���� � �����  �  �         ����	  9 :           }� � t f     ����nd  (�      �     �� ���        ���� � �����  �  �         ����	  < =           �� � y g     �����e  ��      �     �� ���       ���� � �����  �  �         ����	  > ?           �� � ~ h     ����g  �      �     �� ���       ���� � �����  �  �         ����	  @ A           �� � � i     ����Lh  ��   ��  �     �� ���       ���� � �����  �  �         ����	  B C           �� � j     �����i  �   ��  �     �� ���       ���� � �����  �  �         ����	  D E           �� � k     �����j  �   ��  �     �� ���       ���� � �����  �  �         ����	  G H           �� � l     ����*l  �   ��  �     �� ���       ���� �����  �  �         ����	  I J           �� � m     ����tm  p!   ��  �	     �� ���       ���� �����  �  �         ����	  * +           � � hp d     �����a  8�      �      �� ���        ���� � �����  �  �         ����	  , -           � � ou e     ����$c  ��      �     �� ���        ���� � �����  �  �         ����	  . /           � � vz f     ����nd  (�      �     �� ���        ���� � �����  �  �         ����	  0 1           � � } g     �����e  ��      �     �� ���       ���� � �����  �  �         ����	  2 3           � � �� h     ����g  �      �     �� ���       ���� � �����  �  �         ����	  4 5           � � �� i     ����Lh  ��   ��  �     �� ���       ���� � �����  �  �         ����	  7 8           � � �� j     �����i  �   ��  �     �� ���       ���� � �����  �  �         ����	  9 :           � � �� k     �����j  �   ��  �     �� ���       ���� � �����  �  �         ����	  ; <           � � �� l     ����*l  �   ��  �     �� ���       ���� �����  �  �         ����	  = >           � � �� m     ����tm  p!   ��  �	     �� ���       ���� �����  �  �         ����	  ) *           #i #k d     �����a  8�            �� ���        ���� � �����  �  �         ����	  + ,           *n *p e     ����$c  ��           �� ���        ���� � �����  �  �         ����	  - .           1s 1u f     ����nd  (�           �� ���        ���� � �����  �  �         ����	  / 0           8x 8z g     �����e  ��           �� ���       ���� � �����  �  �         ����	  1 2           ?} ? h     ����g  �           �� ���       ���� � �����  �  �         ����	  3 4           F� F� i     ����Lh  ��   ��       �� ���       ���� � �����  �  �         ����	  6 7           M� M� j     �����i  �   ��       �� ���       ���� � �����  �  �         ����	  8 9           T� T� k     �����j  �   ��       �� ���       ���� � �����  �  �         ����	  : ;           [� [� l     ����*l  �   ��       �� ���       ���� �����  �  �         ����	  < =           b� b� m     ����tm  p!   ��  	     �� ���       ���� �����  �  �         ����	    !           � � gn d     �����a  8�            �� ���        ���� � �����  �  �         ����	  " #           � � ns e     ����$c  ��           �� ���        ���� � �����  �  �         ����	  $ %           � � ux f     ����nd  (�           �� ���        ���� � �����  �  �         ����	  & '           � � |} g     �����e  ��           �� ���       ���� � �����  �  �         ����	  ( )           � � �� h     ����g  �           �� ���       ���� � �����  �  �         ����	  * +           � � �� i     ����Lh  ��   ��       �� ���       ���� � �����  �  �         ����	  , -           � � �� j     �����i  �   ��       �� ���       ���� � �����  �  �         ����	  . /           � � �� k     �����j  �   ��       �� ���       ���� � �����  �  �         ����	  0 1           � � �� l     ����*l  �   ��       �� ���       ���� �����  �  �         ����	  2 3           � � �� m     ����tm  p!   ��  	     �� ���       ���� �����  �  �         ����
  6 7           |� v j d     ����J`  x�      A      �� ���        ���� � �����  �  �         ����
  8 9           �� { o e     �����a  �      A     �� ���        ���� � �����  �  �         ����
  : ;           �� � t f     �����b  h�      A     �� ���        ���� � �����  �  �         ����
  = >           �� � y g     ����(d  �      A     �� ���       ���� � �����  �  �         ����
  ? @           �� � ~ h     ����re  X�      A     �� ���       ���� � �����  �  �         ����
  A B           �� � � i     �����f  ��   ��  A     �� ���       ���� � �����  �  �         ����
  C D           �� � j     ����h  H�   ��  A     �� ���       ���� � �����  �  �         ����
  E F           �� � k     ����Pi  ��   ��  A     �� ���       ���� � �����  �  �         ����
  H I           �� � l     �����j  8�   ��  A     �� ���       ���� �����  �  �         ����
  J K           �� � m     �����k  �   ��  A	     �� ���       ���� �����  �  �         ����
  * +           � � up d     ����J`  x�      P      �� ���        ���� � �����  �  �         ����
  , -           � � |u e     �����a  �      P     �� ���        ���� � �����  �  �         ����
  . /           � � �z f     �����b  h�      P     �� ���        ���� � �����  �  �         ����
  0 1           � � � g     ����(d  �      P     �� ���       ���� � �����  �  �         ����
  2 3           � � �� h     ����re  X�      P     �� ���       ���� � �����  �  �         ����
  4 5           � � �� i     �����f  ��   ��  P     �� ���       ���� � �����  �  �         ����
  7 8           � � �� j     ����h  H�   ��  P     �� ���       ���� � �����  �  �         ����
  9 :           � � �� k     ����Pi  ��   ��  P     �� ���       ���� � �����  �  �         ����
  ; <           � �� l     �����j  8�   ��  P     �� ���       ���� �����  �  �         ����
  = >           � 	�� m     �����k  �   ��  P	     �� ���       ���� �����  �  �         ����
  ) *           0i 0k d     ����J`  x�      _      �� ���        ���� � �����  �  �         ����
  + ,           7n 7p e     �����a  �      _     �� ���        ���� � �����  �  �         ����
  - .           >s >u f     �����b  h�      _     �� ���        ���� � �����  �  �         ����
  / 0           Ex Ez g     ����(d  �      _     �� ���       ���� � �����  �  �         ����
  1 2           L} L h     ����re  X�      _     �� ���       ���� � �����  �  �         ����
  3 4           S� S� i     �����f  ��   ��  _     �� ���       ���� � �����  �  �         ����
  6 7           Z� Z� j     ����h  H�   ��  _     �� ���       ���� � �����  �  �         ����
  8 9           a� a� k     ����Pi  ��   ��  _     �� ���       ���� � �����  �  �         ����
  : ;           h� h� l     �����j  8�   ��  _     �� ���       ���� �����  �  �         ����
  < =           o� o� m     �����k  �   ��  _	     �� ���       ���� �����  �  �         ����
    !           � � pw d     ����J`  x�      n      �� ���        ���� � �����  �  �         ����
  " #           � � w| e     �����a  �      n     �� ���        ���� � �����  �  �         ����
  $ %           � � ~� f     �����b  h�      n     �� ���        ���� � �����  �  �         ����
  & '           � � �� g     ����(d  �      n     �� ���       ���� � �����  �  �         ����
  ( )           � � �� h     ����re  X�      n     �� ���       ���� � �����  �  �         ����
  * +           � � �� i     �����f  ��   ��  n     �� ���       ���� � �����  �  �         ����
  , -           � � �� j     ����h  H�   ��  n     �� ���       ���� � �����  �  �         ����
  . /           � � �� k     ����Pi  ��   ��  n     �� ���       ���� � �����  �  �         ����
  0 1           � � �� l     �����j  8�   ��  n     �� ���       ���� �����  �  �         ����
  2 3           � � �� m     �����k  �   ��  n	     �� ���       ���� �����  �  �         ����  7 8           �� v j d     �����U  �      �      �� ���        ���� � �����  �  �         ����  9 :           �� { o e     ����W  `      �     �� ���        ���� � �����  �  �         ����  ; <           �� � t f     ����RX  �#      �     �� ���        ���� � �����  �  �         ����  > ?           �� � y g     �����Y  P3      �     �� ���       ���� � �����  �  �         ����  @ A           �� � ~ h     �����Z  �B      �     �� ���       ���� � �����  �  �         ����  B C           �� � � i     ����0\  @R   ��  �     �� ���       ���� � �����  �  �         ����  D E           �� � j     ����z]  �a   ��  �     �� ���       ���� � �����  �  �         ����  F G           �� � k     �����^  0q   ��  �     �� ���       ���� � �����  �  �         ����  I J           �� � l     ����`  ��   ��  �     �� ���       ���� �����  �  �         ����  K L           �� � m     ����Xa   �   ��  �	     �� ���       ���� �����  �  �         ����  + ,           � � �p d     �����U  �      �      �� ���        ���� � �����  �  �         ����  - .           � � �u e     ����W  `      �     �� ���        ���� � �����  �  �         ����  / 0           � � �z f     ����RX  �#      �     �� ���        ���� � �����  �  �         ����  1 2           � � � g     �����Y  P3      �     �� ���       ���� � �����  �  �         ����  3 4           � � �� h     �����Z  �B      �     �� ���       ���� � �����  �  �         ����  5 6           � � �� i     ����0\  @R   ��  �     �� ���       ���� � �����  �  �         ����  8 9           � �� j     ����z]  �a   ��  �     �� ���       ���� � �����  �  �         ����  : ;           � 
�� k     �����^  0q   ��  �     �� ���       ���� � �����  �  �         ����  < =           � �� l     ����`  ��   ��  �     �� ���       ���� �����  �  �         ����  > ?           � �� m     ����Xa   �   ��  �	     �� ���       ���� �����  �  �         ����  * +           =i =k d     �����U  �      �      �� ���        ���� � �����  �  �         ����  , -           Dn Dp e     ����W  `      �     �� ���        ���� � �����  �  �         ����  . /           Ks Ku f     ����RX  �#      �     �� ���        ���� � �����  �  �         ����  0 1           Rx Rz g     �����Y  P3      �     �� ���       ���� � �����  �  �         ����  2 3           Y} Y h     �����Z  �B      �     �� ���       ���� � �����  �  �         ����  4 5           `� `� i     ����0\  @R   ��  �     �� ���       ���� � �����  �  �         ����  7 8           g� g� j     ����z]  �a   ��  �     �� ���       ���� � �����  �  �         ����  9 :           n� n� k     �����^  0q   ��  �     �� ���       ���� � �����  �  �         ����  ; <           u� u� l     ����`  ��   ��  �     �� ���       ���� �����  �  �         ����  = >           |� |� m     ����Xa   �   ��  �	     �� ���       ���� �����  �  �         ����    !           � � y� d     �����U  �      �      �� ���        ���� � �����  �  �         ����  " #           � � �� e     ����W  `      �     �� ���        ���� � �����  �  �         ����  $ %           � � �� f     ����RX  �#      �     �� ���        ���� � �����  �  �         ����  & '           � � �� g     �����Y  P3      �     �� ���       ���� � �����  �  �         ����  ( )           � � �� h     �����Z  �B      �     �� ���       ���� � �����  �  �         ����  * +           � � �� i     ����0\  @R   ��  �     �� ���       ���� � �����  �  �         ����  , -           � � �� j     ����z]  �a   ��  �     �� ���       ���� � �����  �  �         ����  . /           � � �� k     �����^  0q   ��  �     �� ���       ���� � �����  �  �         ����  0 1           � � �� l     ����`  ��   ��  �     �� ���       ���� �����  �  �         ����  2 3           � �� m     ����Xa   �   ��  �	     �� ���       ���� �����  �  �         ����  8 9           �� v j d     ����jc  ��      �      �� ���        ���� � �����  �  �         ����  : ;           �� { o e     �����d  p�      �     �� ���        ���� � �����  �  �         ����  < =           �� � t f     �����e  ��      �     �� ���        ���� � �����  �  �         ����  ? @           �� � y g     ����Hg  `�      �     �� ���       ���� � �����  �  �         ����  A B           �� � ~ h     �����h  ��      �     �� ���       ���� � �����  �  �         ����  C D           �� � � i     �����i  P�   ��  �     �� ���       ���� � �����  �  �         ����  E F           �� � j     ����&k  �   ��  �     �� ���       ���� � �����  �  �         ����  G H           �� � k     ����pl  @   ��  �     �� ���       ���� � �����  �  �         ����  J K           �� � l     �����m  �$   ��  �     �� ���       ���� �����  �  �         ����  L M           �� � m     ����o  04   ��  �	     �� ���       ���� �����  �  �         ����  + ,           � � �p d     ����jc  ��            �� ���        ���� � �����  �  �         ����  - .           � � �u e     �����d  p�           �� ���        ���� � �����  �  �         ����  / 0           � � �z f     �����e  ��           �� ���        ���� � �����  �  �         ����  1 2           � � � g     ����Hg  `�           �� ���       ���� � �����  �  �         ����  3 4           � �� h     �����h  ��           �� ���       ���� � �����  �  �         ����  5 6           � �� i     �����i  P�   ��       �� ���       ���� � �����  �  �         ����  8 9           � �� j     ����&k  �   ��       �� ���       ���� � �����  �  �         ����  : ;           � �� k     ����pl  @   ��       �� ���       ���� � �����  �  �         ����  < =           � �� l     �����m  �$   ��       �� ���       ���� �����  �  �         ����  > ?           � #�� m     ����o  04   ��  	     �� ���       ���� �����  �  �         ����  * +           Ji Jk d     ����jc  ��            �� ���        ���� � �����  �  �         ����  , -           Qn Qp e     �����d  p�           �� ���        ���� � �����  �  �         ����  . /           Xs Xu f     �����e  ��           �� ���        ���� � �����  �  �         ����  0 1           _x _z g     ����Hg  `�           �� ���       ���� � �����  �  �         ����  2 3           f} f h     �����h  ��           �� ���       ���� � �����  �  �         ����  4 5           m� m� i     �����i  P�   ��       �� ���       ���� � �����  �  �         ����  7 8           t� t� j     ����&k  �   ��       �� ���       ���� � �����  �  �         ����  9 :           {� {� k     ����pl  @   ��       �� ���       ���� � �����  �  �         ����  ; <           �� �� l     �����m  �$   ��       �� ���       ���� �����  �  �         ����  = >           �� �� m     ����o  04   ��  	     �� ���       ���� �����  �  �         ����    !           � � �� d     ����jc  ��      "      �� ���        ���� � �����  �  �         ����  " #           � � �� e     �����d  p�      "     �� ���        ���� � �����  �  �         ����  $ %           � � �� f     �����e  ��      "     �� ���        ���� � �����  �  �         ����  & '           � � �� g     ����Hg  `�      "     �� ���       ���� � �����  �  �         ����  ( )           � � �� h     �����h  ��      "     �� ���       ���� � �����  �  �         ����  * +           � � �� i     �����i  P�   ��  "     �� ���       ���� � �����  �  �         ����  , -           � � �� j     ����&k  �   ��  "     �� ���       ���� � �����  �  �         ����  . /           � �� k     ����pl  @   ��  "     �� ���       ���� � �����  �  �         ����  0 1           � �� l     �����m  �$   ��  "     �� ���       ���� �����  �  �         ����  2 3           � �� m     ����o  04   ��  "	     �� ���       ���� �����  �  �         ����  8 9           �� v j d     �����d  ��      O      �� ���        ���� � �����  �  �         ����  : ;           �� { o e     ����Df  0�      O     �� ���        ���� � �����  �  �         ����  < =           �� � t f     �����g  ��      O     �� ���        ���� � �����  �  �         ����  ? @           �� � y g     �����h   �      O     �� ���       ���� � �����  �  �         ����  A B           �� � ~ h     ����"j  ��      O     �� ���       ���� � �����  �  �         ����  C D           �� � � i     ����lk  	   ��  O     �� ���       ���� � �����  �  �         ����  E F           �� � j     �����l  �   ��  O     �� ���       ���� � �����  �  �         ����  G H           �� � k     ���� n   (   ��  O     �� ���       ���� � �����  �  �         ����  J K           �� � l     ����Jo  x7   ��  O     �� ���       ���� �����  �  �         ����  L M           �� � m     �����p  �F   ��  O	     �� ���       ���� �����  �  �         ����  + ,           � � �p d     �����d  ��      ^      �� ���        ���� � �����  �  �         ����  - .           � � �u e     ����Df  0�      ^     �� ���        ���� � �����  �  �         ����  / 0           � � �z f     �����g  ��      ^     �� ���        ���� � �����  �  �         ����  1 2           � � g     �����h   �      ^     �� ���       ���� � �����  �  �         ����  3 4           � �� h     ����"j  ��      ^     �� ���       ���� � �����  �  �         ����  5 6           � �� i     ����lk  	   ��  ^     �� ���       ���� � �����  �  �         ����  8 9           � �� j     �����l  �   ��  ^     �� ���       ���� � �����  �  �         ����  : ;           � �� k     ���� n   (   ��  ^     �� ���       ���� � �����  �  �         ����  < =           �  �� l     ����Jo  x7   ��  ^     �� ���       ���� �����  �  �         ����  > ?           � &�� m     �����p  �F   ��  ^	     �� ���       ���� �����  �  �         ����  * +           Mi Mk d     �����d  ��      m      �� ���        ���� � �����  �  �         ����  , -           Tn Tp e     ����Df  0�      m     �� ���        ���� � �����  �  �         ����  . /           [s [u f     �����g  ��      m     �� ���        ���� � �����  �  �         ����  0 1           bx bz g     �����h   �      m     �� ���       ���� � �����  �  �         ����  2 3           i} i h     ����"j  ��      m     �� ���       ���� � �����  �  �         ����  4 5           p� p� i     ����lk  	   ��  m     �� ���       ���� � �����  �  �         ����  7 8           w� w� j     �����l  �   ��  m     �� ���       ���� � �����  �  �         ����  9 :           ~� ~� k     ���� n   (   ��  m     �� ���       ���� � �����  �  �         ����  ; <           �� �� l     ����Jo  x7   ��  m     �� ���       ���� �����  �  �         ����  = >           �� �� m     �����p  �F   ��  m	     �� ���       ���� �����  �  �         ����    !           � � �� d     �����d  ��      |      �� ���        ���� � �����  �  �         ����  " #           � � �� e     ����Df  0�      |     �� ���        ���� � �����  �  �         ����  $ %           � � �� f     �����g  ��      |     �� ���        ���� � �����  �  �         ����  & '           � � �� g     �����h   �      |     �� ���       ���� � �����  �  �         ����  ( )           � � �� h     ����"j  ��      |     �� ���       ���� � �����  �  �         ����  * +           � � �� i     ����lk  	   ��  |     �� ���       ���� � �����  �  �         ����  , -           � � �� j     �����l  �   ��  |     �� ���       ���� � �����  �  �         ����  . /           � �� k     ���� n   (   ��  |     �� ���       ���� � �����  �  �         ����  0 1           � �� l     ����Jo  x7   ��  |     �� ���       ���� �����  �  �         ����  2 3           � �� m     �����p  �F   ��  |	     �� ���       ���� �����  �  �          ����                       2   `	  �       �      �   �        ���� � �������������          ����               $        0   ~	  �       �     �   �        ���� � �������������          ����               )        1   �	  8       �     �   �        ���� � �������������          ����  	 
            .        1   �	  t       �     �   �       ���� � �������������          ����              " 3 !       2   �	  �       �     �   �       ���� � �������������          ����              % 8 #       3   �	  �       �     �   �       ���� � �������������          ����              ( = %       3   
  (       �     �   �       ���� � �������������          ����             ! + B '       4   2
  d       �     �   �       ���� � �������������          ����             # . G )       4   P
  �       �     �   �       ���� � �������������          ����             % 1 L +       5   n
  �       �	     �   �       ���� � �������������          ����               :        S   �
  �        �      �   �        ���� � �������������          ����   	           ! ?        U   "  f!       �     �   �        ���� � �������������          ����  
            $ D        W   ^  "       �     �   �        ���� � �������������          ����              ' I        Y   �  �"       �     �   �       ���� � �������������          ����              * N         Z   �  �#       �     �   �       ���� � �������������          ����             ! - S "       \     6$       �     �   �       ���� � �������������          ����             $ 0 X $       ^   N  �$       �     �   �       ���� � �������������          ����             ' 3 ] &       `   �  �%       �     �   �       ���� � �������������          ����             * 6 b (       b   �  R&       �     �   �       ���� � �������������          ����             - 9 g *       c     '       �	     �   �       ���� � �������������         ����  	 
           % T        �   �  �7       �      �   �        ���� � �������������         ����              ) Y        �   L  09       �     �   �        ���� � �������������         ����               - ^        �   �  �:       �     �   �        ���� � �������������         ����             # 1 c        �       <       �     �   �       ���� � �������������         ����             & 5 h "       �   Z  h=       �     �   �       ���� � �������������         ����             ) 9 m %       �   �  �>       �     �   �       ���� � �������������         ����             , = r (       �     8@       �     �   �       ���� � �������������         ����             / A w +       �   h  �A       �     �   �       ���� � �������������         ����             2 E | .       �   �  C       �     �   �       ���� � �������������         ����             5 I � 1       �     pD       �	     �   �       ���� � �������������         ����             " 6 m        �   �  �\       �      �   �        ���� � �������������         ����             % : s !       �   �  �^       �     �   �        ���� � �������������         ����             ( > y $       �   t  Da       �     �   �        ���� � �������������         ����             + B  '       �   �  �c       �     �   �       ���� � �������������         ����             . F � *         d  �e       �     �   �       ���� � �������������         ����             1 J � -         �  Lh       �     �   �       ���� � �������������         ����             4 N � 0         T  �j       �     �   �       ���� � �������������         ����             7 R � 3         �  �l       �     �   �       ���� � �������������         ����             : V � 6         D  To       �     �   �       ���� � �������������         ����             = Z � 9       #  �  �q       �	     �   �       ���� � �������������         ����             ) F � %       z  �  ��       �      �   �        ���� � �������������         ����             , J � (       �  2  ,�       �     �   �        ���� � �������������         ����             / N � +       �  �  ��       �     �   �        ���� � �������������         ����             2 R � .       �  ^  4�       �     �   �       ���� � �������������         ����             5 V � 1       �  �  ��       �     �   �       ���� � �������������         ����             8 Z � 4       �  �  <�       �     �   �       ���� � �������������         ����             ; ^ � 7       �     ��       �     �   �       ���� � �������������         ����             > b � :       �  �  D�       �     �   �       ���� � �������������         ����              A f � =       �  L  ȯ    
   �     �   �       ���� � �������������         ����  ! "          D j � @       �  �  L�    	   �	     �   �       ���� � �������������         ����             0 U � ,       A  :   ��       �      �   �        ���� � �������������         ����             4 Y � /       N  �   ��       �     �   �        ���� � �������������         ����             8 ] � 2       Z  �!  n�       �     �   �        ���� � �������������         ����             < a � 5       g  V"  Z�       �     �   �       ���� � �������������         ����             @ e � 8       s  
#  F�       �     �   �       ���� � �������������         ����             D i � ;       �  �#  2�       �     �   �       ���� � �������������         ����             H m � >       �  r$  �       �     �   �       ���� � �������������         ����    !          L q � A       �  &%  
   	   �     �   �       ���� � �������������         ����  " #          P u � D       �  �%  �      �     �   �       ���� � �������������         ����  $ %          T y � G       �  �&  �      �	     �   �       ���� � �������������         ����             @ d � 2       O  ^)  �J      �      �   �        ���� � �����  �  �         ����             D i � 6       `  0*  �Q      �     �   �        ���� � �����  �  �         ����             H n � :       p  +  X      �     �   �        ���� � �����  �  �         ����             L s � >       �  �+  �^      �     �   �       ���� � �����  �  �         ����             P x � B       �  �,  0e      �     �   �       ���� � �����  �  �         ����              T } � F       �  x-  �k   	   �     �   �       ���� � �����  �  �         ����  ! "          X � � J       �  J.  Pr      �     �   �       ���� � �����  �  �         ����  # $          \ � � N       �  /  �x      �     �   �       ���� � �����  �  �         ����  % &          ` � R       �  �/  p      �     �   �       ���� � �����  �  �         ����  ' (          d � V       �  �0   �      �	     �   �       ���� � �����  �  �         ����             P | � B       �  4  H�      �      �   �        ���� � �����  �  �         ����             T � � F       �  �4  ��      �     �   �        ���� � �����  �  �         ����             X �  J       �  �5  (�      �     �   �        ���� � �����  �  �         ����             \ � N       �  �6  ��   	   �     �   �       ���� � �����  �  �         ����    !          ` � R         �7  �      �     �   �       ���� � �����  �  �         ����  " #          d � V         �8  x�      �     �   �       ���� � �����  �  �         ����  $ %          h � Z       0  �9  �      �     �   �       ���� � �����  �  �         ����  & '          l � #^       F  �:  X      �     �   �       ���� � �����  �  �         ����  ( )          p � *b       [  �;  �      �     �   �       ���� � �����  �  �         ����  * +          t � 1f       q  x<  8       �	     �   �       ���� � -  �  �  �         ����             _ � Q       l  8@  0�      �      �   �        ����	 � �����  �  �         ����             c � "U       �  FA  ��   
   �     �   �        ����	 � �����  �  �         ����              g � )Y       �  TB  H�      �     �   �        ����	 � �����  �  �         ����  ! "          k � 0]       �  bC  ԡ      �     �   �       ����	 � �����  �  �         ����  # $          o � 7a       �  pD  `�      �     �   �       ����	 � �����  �  �         ����  % &          s � >e       �  ~E  �      �     �   �       ����	 � �����  �  �         ����  ' (          w � Ei         �F  x�      �     �   �       ����	 � �����  �  �         ����  ) *          { � Lm       )  �G  �      �     �   �       ����	 � �����  �  �         ����  + ,           � Sq       D  �H  ��       �     �   �       ����	 � �����  �  �         ����  - .          � � Zu       _  �I  �   ��  �	     �   �       ����	 � 7  �  �  �         ����             n � C`       �  �M  :Y   	   �      �   �        ����
 � �����  �  �         ����    !          s � Jd       �  O  f      �     �   �        ����
 � �����  �  �         ����  " #          x � Qh       �  FP  s      �     �   �        ����
 � �����  �  �         ����  $ %          } � Xl       �  rQ  �      �     �   �       ����
 � �����  �  �         ����  & '          � � _p       	  �R  ʌ      �     �   �       ����
 � �����  �  �         ����  ( )          � � ft       7	  �S  ��      �     �   �       ����
 � �����  �  �         ����  * +          � � mx       X	  �T  ��      �     �   �       ����
 � �����  �  �         ����  , -          � � t|       y	  "V  v�   ��  �     �   �       ����
 � �����  �  �         ����  . /          � � {�       �	  NW  Z�   ��  �     �   �       ����
 � �����  �  �         ����  0 1          � � ��       �	  zX  >�   ��  �	     �   �       ����
 7  �  �  �         ����  ! "          � � jn d     .  *]  �]      �      �   �        ���� � �����  �  �         ����  # $          � � qs e     U  t^  pm      �     �   �        ���� � �����  �  �         ����  % &          � � xx f     }  �_  �|      �     �   �        ���� � �����  �  �         ����  ' (          � � } g     �  a  `�      �     �   �       ���� � �����  �  �         ����  ) *          � � �� h     �  Rb  ؛      �     �   �       ���� � �����  �  �         ����  + ,          � � �� i     �  �c  P�   ��  �     �   �       ���� � �����  �  �         ����  - .          � � �� j       �d  Ⱥ   ��  �     �   �       ���� � �����  �  �         ����  / 0          � � �� k     C  0f  @�   ��  �     �   �       ���� � �����  �  �         ����  1 2          � � �� l     j  zg  ��   ��  �     �   �       ���� �����  �  �         ����  3 4          � � �� m     �  �h  0�   ��  �	     �   �       ���� A  �  �  �            ��A�+�2    %� � d     i  ĸ  E                 �    ������� � �����  �  �            ��X�E�2    -�� � e     �  ��  �d                �    ������� � �����  �  �            ��o�_�2    5�� � f        ��  Ą                �    ������� � �����  �  �            ���y2    =�� g     ]   d�  ��                �   ������� � �����  �  �            ���(�(2    E�
� h     �   D�  ��                �   ������� � �����  �  �            ���@�C2    M�i     !  $�  d�   ��            �   ������� � �����  �  �            ���X�^2    U�
j     R!  �  D   ��            �   ������� � �����  �  �            ���p�y2    ]�k     �!  ��  $$   ��            �   ������� � �����  �  �            ������2    e�"l     �!  ��  D   ��            �   �������  �����  �  �            ����2    m�(m     G"  ��  �c   ��   	         �   ������� 	   �  �  �            ���,�X2    4�� � d     �  ��  �T      '       %   �    ������� � �����  �  �            ���I�o2    <�� � e     �  ��  �t      '      %   �    ������� � �����  �  �            ���f��2    D�� � f     5   t�  ��      '      %   �    ������� � �����  �  �            �����2    L�� g     �   T�  ��      '      %   �   ������� � �����  �  �            ����2    T�
� h     �   4�  t�      '      %   �   ������� � �����  �  �            ��1�0�2    \�i     )!  �  T�   ��  '      %   �   ������� � �����  �  �            ��M�E�2    d�
j     {!  ��  4   ��  '      %   �   ������� � �����  �  �            ��i�Z�2    l�k     �!  ��  4   ��  '      %   �   ������� � �����  �  �            ���o2    t�"l     "  ��  �S   ��  '      %   �   �������  �����  �  �            ���1�'2    |�(m     p"  ��  �s   ��  ' 	     %   �   ������� 	G   �  �  �            ���L�L2    �� �� d     s   �   I      ;       9   �    ������� � �����  �  �            ���f�f2    � �� e     �  �  �h      ;      9   �    ������� � �����  �  �            ������2    ��� f        ��  ��      ;      9   �    ������� � �����  �  �            ����2    �� g     h   ��  ��      ;      9   �   ������� � �����  �  �            ����2    h     �   ��  ��      ;      9   �   ������� � �����  �  �            ��8�8�2    i     !  `�  `�   ��  ;      9   �   ������� � �����  �  �            ��Q�Q�2    j     \!  @�  @   ��  ;      9   �   ������� � �����  �  �            ��jj2    $k     �!   �   (   ��  ;      9   �   ������� � �����  �  �            ����2    &*&l      "   �   H   ��  ;      9   �   �������  �����  �  �            ���6�62    .0.$m     Q"  ��  �g   ��  ; 	     9   �   ������� 	y   �  �  �            ��+�A�2    /�� � d     �  x�  �P      Q       N   �    ������� � �����  �  �            ��E�X�2    7�� � e     �  X�  �p      Q      N   �    ������� � �����  �  �            ��_�o�2    ?�� � f     *   8�  ��      Q      N   �    ������� � �����  �  �            ��y�2    G�� g     |   �  ��      Q      N   �   ������� � �����  �  �            ���(�(2    O�
� h     �   ��  x�      Q      N   �   ������� � �����  �  �            ���C�@2    W�i     !  ��  X�   ��  Q      N   �   ������� � �����  �  �            ���^�X2    _�
j     q!  ��  8   ��  Q      N   �   ������� � �����  �  �            ���y�p2    g�k     �!  ��  0   ��  Q      N   �   ������� � �����  �  �            ������2    o�"l     "  x�  �O   ��  Q      N   �   �������  �����  �  �            ����2    w�(m     f"  X�  �o   ��  Q 	     N   �   ������� 	�   �  �  �            ���X�,2    a*� d     ^  ��  A      g       c   �    ������� � �����  �  �            ���o�I2    h2� e     �  h�  �`      g      c   �    ������� � �����  �  �            �����f2    o:� f        H�  Ȁ      g      c   �    ������� � �����  �  �            �����2    vB� g     S   (�  ��      g      c   �   ������� � �����  �  �            ����2    %}Jh     �   �  ��      g      c   �   ������� � �����  �  �            ��0�1�2    +�R
i     �   ��  h�   ��  g      c   �   ������� � �����  �  �            ��E�M�2    1�Zj     H!  ��  H    ��  g      c   �   ������� � �����  �  �            ��Z�i�2    7�bk     �!  ��  (    ��  g      c   �   ������� � �����  �  �            ��o�2    =�jl     �!  ��  @   ��  g      c   �   �������  �����  �  �            ���'�12    C�r"m     ="  h�  �_   ��  g 	     c   �   ������� 	�   �  �  �             t�t�
2    �� �� d     }  <�  �L      �       {   �    ������� � �����  �  �             ��
2    � �� e     �  �  �l      �      {   �    ������� � �����  �  �             �-�-
2    ��� f         ��  ��      �      {   �    ������� � �����  �  �             �F�F
2    �� g     r   ܾ  ��      �      {   �   ������� � �����  �  �             �_�_
2    h     �   ��  |�      �      {   �   ������� � �����  �  �             �x�x
2    i     !  ��  \�   ��  �      {   �   ������� � �����  �  �             ��
2    j     g!  |�  <   ��  �      {   �   ������� � �����  �  �             ��
2    $k     �!  \�  ,   ��  �      {   �   ������� � �����  �  �             4�4�
2    $*&l     
"  <�  �K   ��  �      {   �   �������  �����  �  �             L�L�
2    ,0.$m     ["  �  �k   ��  � 	     {   �   ������� 	  �  �  �         ����   # $            d �         	      �        a        ���        ����c   �������������         ����   % &            g �            >  |        a       ���        ����c   �������������         ����   ' (            j �            \  �        a       ���        ����c   �������������         ����   ) *            m �            z  �        a       ���       ����c   �������������         ����   + ,            p �            �  0        a       ���       ����c   �������������         ����   - .            s �            �  l        a       ���       ����c   �������������         ����   / 0            v �            �  �        a       ���       ����c   �������������         ����   1 2            y �            �  �        a       ���       ����c   �������������         ����   3 4            | �                       a       ���       ����c   �������������         ����   5 6             �            .  \        a	       ���       ����c   �������������         ����  " #            d �            ,  h        �        ���        ����c   �������������         ����  $ %            g �            J  �        �       ���        ����c   �������������         ����  & '            j �            h  �        �       ���        ����c   �������������         ����  ( )            m �            �          �       ���       ����c   �������������         ����  * +            p �            �  H        �       ���       ����c   �������������         ����  , -            s �         	   �  �        �       ���       ����c   �������������         ����  . /            v �         	   �  �        �       ���       ����c   �������������         ����  0 1            y �         
   �  �        �       ���       ����c   �������������         ����  2 3            | �         
     8        �       ���       ����c   �������������         ����  4 5             �            :  t        �	       ���       ����c   �������������         ����  ! #            d �            �   �         2        ���        ����c   �������������         ����  # %            g �            �   �        2       ���        ����c   �������������         ����  % '            j �                      2       ���        ����c   �������������         ����  ' )            m �            "  D        2       ���       ����c   �������������         ����  ) +            p �            @  �        2       ���       ����c   �������������         ����  + -            s �            ^  �        2       ���       ����c   �������������         ����  - /            v �            |  �        2       ���       ����c   �������������         ����  / 1            y �            �  4        2       ���       ����c   �������������         ����  1 3            | �            �  p        2       ���       ����c   �������������         ����  3 5             �         	   �  �        2	       ���       ����c   �������������         ����  " #            d �         !   �  /        �        ���        ����c   �������������         ����  $ %            g �         (   �  �        �       ���        ����c   �������������         ����  & '            j �         )             �       ���        ����c   �������������         ����  ( )            m �         )   *  T        �       ���       ����c   �������������         ����  * +            p �         *   H  �        �       ���       ����c   �������������         ����  , -            s �         +   f  �        �       ���       ����c   �������������         ����  . /            v �         +   �          �       ���       ����c   �������������         ����  0 1            y �         ,   �  D        �       ���       ����c   �������������         ����  2 3            | �         ,   �  �        �       ���       ����c   �������������         ����  4 5             �         -   �  �        �	       ���       ����c   �������������         ����  # $            d �            @  �        �        ���        ����c   �������������         ����  % &            g �             ^  �        �       ���        ����c   �������������         ����  ' (            j �         !   |  �        �       ���        ����c   �������������         ����  ) *            m �         !   �  4        �       ���       ����c   �������������         ����  + ,            p �         "   �  p        �       ���       ����c   �������������         ����  - .            s �         #   �  �        �       ���       ����c   �������������         ����  / 0            v �         #   �  �        �       ���       ����c   �������������         ����  1 2            y �         $     $        �       ���       ����c   �������������         ����  3 4            | �         $   0  `        �       ���       ����c   �������������         ����  5 6             �         %   N  �        �	       ���       ����c   �������������         ����  " #            d �            �  F        d        ���        ����c   �������������         ����  $ %            g �            �  �	        d       ���        ����c   �������������         ����  & '            j �            �  �	        d       ���        ����c   �������������         ����  ( )            m �            
  
        d       ���       ����c   �������������         ����  * +            p �            (  P
        d       ���       ����c   �������������         ����  , -            s �            F  �
        d       ���       ����c   �������������         ����  . /            v �            d  �
        d       ���       ����c   �������������         ����  0 1            y �            �          d       ���       ����c   �������������         ����  2 3            | �            �  @        d       ���       ����c   �������������         ����  4 5             �            �  |        d	       ���       ����c   �������������                  2                   �  �    $   �       �   �    ������ � �������������                  2                         #   �      �   �    ������ � �������������                  2                      @    !   �      �   �    ������ � �������������               
  	 2                    >  |        �      �   �   ������ � �������������              
  	  2    $               \  �       �      �   �   ������ � �������������                  2    (               z  �       �      �   �   ������ � �������������                  2    ,               �  0       �      �   �   ������ � �������������                  2    0               �  l       �      �   �   ������ � �������������                  2    4               �  �       �      �   �   ������ � �������������                  2    8               �  �       � 	     �   �   ������ � �������������                  2    % #           !   j  >    "   �       �   �    ������� � �������������                  2    ) (           #   �  �    !   �      �   �    ������� � �������������                  2    - -           %   �  �       �      �   �    ������� � �������������                   2    1 2           '     Z       �      �   �   ������� � �������������              ! $   2    5 7           )   Z         �      �   �   ������� � �������������              % (  " 2    9 <           *   �  �       �      �   �   ������� � �������������              ) , " % 2    = A           ,   �  v       �      �   �   ������� � �������������              - 0 % ( 2    A F           .     *       �      �   �   ������� � �������������              1 4 ( + 2    E K           0   J  �       �      �   �   ������� � �������������              5 8 + . 2    I P           2   �  �       � 	     �   �   ������� � �������������              . 2 # ' 2    6 >          L   v  �        �       �   �    ������� � �������������              3 8 ' , 2    : C !         P   �  @       �      �   �    ������� � �������������              8 > + 1 2    > H $         S   *  �        �      �   �    ������� � �������������              = D / 6 2    B M '         W   �  "       �      �   �   ������� � �������������              B J 3 ; 2    F R *         Z   �  x#       �      �   �   ������� � �������������              G P 7 @ 2    J W -         ^   8	  �$       �      �   �   ������� � �������������              L V ; E 2    N \ 0         b   �	  H&       �      �   �   ������� � �������������              Q \ ? J 2    R a 3         e   �	  �'       �      �   �   ������� � �������������              V b C O 2    V f 6         i   F
  )       �      �   �   ������� � �������������              [ h G T 2    Z k 9         l   �
  �*       � 	     �   �   ������� � �������������              O _ : J 2    F X &        �     (<       �       �        ˹I���� � �������������              V g @ P 2    J ] )        �   �  �>       �      �        ˹I���� � �������������              ] o F V 2    N b ,         �   �  �@       �      �        ˹I���� � �������������              d w L \ 2    R g / #       �   p  0C       �      �       ˹I���� � �������������              k  R b 2    V l 2 &       �   �  �E       �      �       ˹I���� � �������������              r � X h 2    Z q 5 )       �   `  �G       �      �       ˹I���� � �������������              y � ^ n 2    ^ v 8 ,       �   �  8J       �      �       ˹I���� � �������������              � � d t 2    b { ; /       �   P  �L       �      �       ˹I���� � �������������              � � j z 2    f � > 2       �   �  �N       �      �       ˹I���� � �������������              � � p � 2    j � A 5       �   @  @Q       � 	     �       ˹I���� � �������������              ~ � _ q 2    U q - !            �l       �       �       ������ � �������������              � � f y 2    Z v 0 $         �  Dp       �      �       ������ � �������������              � � m � 2    _ { 3 '       (  L  �s       �      �       ������ � �������������              � � t � 2    d � 6 *       1  �  Lw       �      �      ������ � �������������              � � { � 2    i � 9 -       :  x  �z       �      �      ������ � �������������              � � � � 2    n � < 0       C    T~       �      �      ������ � �������������              � � � � 2    s � ? 3       L  �  ؁       �      �      ������ � �������������              � � � � 2    x � B 6       U  :  \�       �      �      ������ � �������������              � � � � 2    } � E 9       ^  �  ��       �      �      ������ � �������������              � � � � 2    � � H <       g  f  d�       � 	     �      ������ � �������������              � � � � 2    m � 4 (       �  �  2�       �       �       j����� � �������������              � � � � 2    r � 7 +       �  r  �       �      �       j����� � �������������              � � � � 2    w � : .       �  &  
�       �      �       j����� � �������������              � � � � 2    | � = 1       �  �  ��       �      �      j����� � �������������              � � � 2    � � @ 4       �  �  ��       �      �      j����� � �������������              � � � 2    � � C 7         B  ��       �      �      j����� � �������������              � � � 2    � � F :         �  ��       �      �      j����� � �������������              '� � 2    � � I =       %  �  ��       �      �      j����� � �������������              2� � 2    � � L @       2  ^  ��       �      �      j����� � �������������              =� � 2    � � O C       >     ~�       � 	     �      j����� � �������������              � (� � 2    � � : .       �  �"        �       �       ϕ����� � �����  �  �              
5� � 2    � � > 2       �  �#  �      �      �       ϕ����� � �����  �  �              B� � 2    � � B 6       �  �$  0$      �      �       ϕ����� � �����  �  �              "O� � 2    � � F :       �  X%  �*      �      �      ϕ����� � �����  �  �              .\� 	2    � � J >         *&  P1      �      �      ϕ����� � �����  �  �              :i� 2    � � N B         �&  �7      �      �      ϕ����� � �����  �  �              Fv� 2    � � R F       /  �'  p>      �      �      ϕ����� � �����  �  �              R�� '2    � � V J       @  �(   E      �      �      ϕ����� � �����  �  �              ^�12    � � Z N       P  r)  �K      �      �      ϕ����� � �����  �  �              j�;2    � � ^ R       a  D*   R      � 	     �      ϕ����� � �����  �  �              N��  2    � � J >         �-  �      �       �       ������ � �����  �  �              \�� ,2    � � N B       /  |.  \�      �      �       ������ � �����  �  �              j�	82    � � R F       D  l/  ̪      �      �       ������ � �����  �  �              x�D2    � � V J       Z  \0  <�      �      �      ������ � �����  �  �              ��P2    � � Z N       o  L1  ��      �      �      ������ � �����  �  �              ��*\2    � � ^ R       �  <2  �      �      �      ������ � �����  �  �              ��5h2    � � b V       �  ,3  ��      �      �      ������ � �����  �  �              ��@t2    � � f Z       �  4  ��      �      �      ������ � �����  �  �              ��K�2    � � j ^       �  5  l�      �      �      ������ � �����  �  �              �V�2    � n b       �  �5  ��   
   � 	     �      ������ � �����  �  �             ��3m2    � � Y M       �  �9  XA      �       �       �������	 � �����  �  �             ��?z2    � � ] Q       �  �:  �K      �      �       �������	 � �����  �  �             �K�2    � � a U       �  �;  pV      �      �       �������	 � �����  �  �             �W�2    � � e Y         �<  �`      �      �      �������	 � �����  �  �             �&c�2    � i ]       2  �=  �k      �      �      �������	 � �����  �  �             �6o�2    � 	m a       M  ?  v      �      �      �������	 � �����  �  �             F{�2    � q e       h  @  ��      �      �      �������	 � �����  �  �             V��2    � u i       �  A  ,�      �      �      �������	 � �����  �  �             $f��2    � y m       �  ,B  ��   	   �      �      �������	 � �����  �  �             3v��2    � !} q       �  :C  D�      � 	     �      �������	 � �����  �  �             Vx�2    � 
h \       �  rG  �      �       �       �������
 � �����  �  �              h��2    � l `       �  �H  �      �      �       �������
 � �����  �  �             1z��2    � p d         �I  �+      �      �       �������
 � �����  �  �             B���2    � t h       >  �J  �8      �      �      �������
 � �����  �  �             S���2    � &x l       _  "L  vE      �      �      �������
 � �����  �  �             d��2    � -| p       �  NM  ZR      �      �      �������
 � �����  �  �             u��2    � 4� t       �  zN  >_   
   �      �      �������
 � �����  �  �             ���!2    � ;� x       �  �O  "l   	   �      �      �������
 � �����  �  �             ���/2     B� |       �  �P  y      �      �      �������
 � �����  �  �             ���=2    I� �       	  �Q  �      � 	     �      �������
 � �����  �  �             ���2    � 2v j       f
  �V  (      �       �       ������� � �����  �  �             ���%2    � 9{ o       �
  �W  �      �      �       ������� � �����  �  �             ���52    � @� t       �
  BY  /      �      �       ������� � �����  �  �             ��E2     G� y       �
  �Z  �>      �      �      ������� � �����  �  �             �$U2    N� ~         �[  N      �      �      ������� � �����  �  �             �8e2    U� �       ,   ]  �]   	   �      �      ������� � �����  �  �             �L%u2    \� �       T  j^  �l      �      �      ������� � �����  �  �             `4�2    c� �       |  �_  p|      �      �      ������� � �����  �  �             tC�2    j� �       �  �`  �      �      �      ������� � �����  �  �             +�R�2    $q� �       �  Hb  `�      � 	     �      ������� � �����  �  �             �a"z2    Y� �       r  pg  �@      �       �       ������� � �����  �  �             v2�2    `� �       �  �h  �R      �      �       ������� � �����  �  �             '�B�2    g� �       �  @j  @e      �      �       ������� � �����  �  �             ;�R�2    n� �       �  �k  �w   
   �      �      ������� � �����  �  �             O�b�2    #u� �       -  m  Љ   	   �      �      ������� � �����  �  �             c�r�2    )|� �       \  xn  �      �      �      ������� � �����  �  �             w���2    /�� �       �  �o  `�      �      �      ������� � �����  �  �             ����2    5�� �       �  Hq  ��      �      �      ������� � �����  �  �             �	�2    ;�� �       �  �r  ��      �      �      ������� � �����  �  �             ��2    A�� �         t  8�      � 	     �      ������� �    �  �  �             ��}�2    '� �       
  �y  �      �       �   	    ioe���� � �����  �  �             �	��2    .�� �       A  >{  d�      �      �   	    ioe���� � �����  �  �             � �	2    5�� �       w  �|  ��   	   �      �   	    ioe���� � �����  �  �             �7�2    <�� �       �  J~  �      �      �   	   ioe���� � �����  �  �             �N�/2    C�� �       �  �  `�      �      �   	   ioe���� � �����  �  �             �e�B2    J�� �         V�  �      �      �   	   ioe���� � �����  �  �             |�U2    Q�� �       R  ܂  (      �      �   	   ioe���� � �����  �  �             ��h2    X�� �       �  b�  \=      �      �   	   ioe���� � �����  �  �             2�{2    _�� �       �  �  �R      �      �   	   ioe���� � �����  �  �             H��2    f�� �       �  n�  h       � 	     �   	   ioe���� �    �  �  �             ��[2    M�� �       :  ��  �J   
   �       �   
    ������ � �����  �  �             ,��o2    T�� �       y  *�  vc   	   �      �   
    ������ � �����  �  �             D��2    [�� �       �  ΐ  |      �      �   
    ������ � �����  �  �             \� �2    b�� �       �  r�  ��      �      �   
   ������ � �����  �  �             t�3�2    i�� �       6  �  J�      �      �   
   ������ � �����  �  �             �F�2    p�� �       u  ��  ��      �      �   
   ������ � �����  �  �             �(Y�2    w�� �       �  ^�  ��      �      �   
   ������ � �����  �  �             �Al�2    ~�� �       �  �  �      �      �   
   ������ � �����  �  �             �Z�2    ��� �       2  ��  �	   ��  �      �   
   ������ � �����  �  �             �s�2    ��� �       q  J�  V(	   ��  � 	     �   
   ������ �    �  �  �             �@U�2    r�� �         ڢ  �-
      �       �       :������ � �����  �  �             �[i�2    y�� �       V  ��  �I
      �      �       :������ � �����  �  �             �v}2    ��� �       �  ^�  �e
      �      �       :������ � �����  �  �             ���2    ��� �       �   �   �
      �      �      :������ � �����  �  �             ��+2    ��� �       .  �   �
      �      �      :������ � �����  �  �             1��@2    ��� �       v  ��  @�
      �      �      :������ � �����  �  �             J��U2    �� �       �  f�  `�
       �      �      :������ � �����  �  �             c��j2    �� �         (�  ��
   ��  �      �      :������ � �����  �  �             |�2    ��       N  �  �   ��  �      �      :������ � �����  �  �             �3	�2    ��       �  ��  �*   ��  � 	     �      :������    �  �  �           ��q  
  
   d                �   �   �        �       �� ��        ������  ����������������         ��q  B D B D  �    t x           �   T  �        �       �� ��        ������  ����������������         ��q  z | z |  �    � �          �              �       �� ��        ������  ����������������         ��q  � � � �  �    � � 6        �     n        �       �� ��        ������  ����������������         ��q  � � � �  �    � � ; ;       �   ~  �        �       �� ��        ������  ����������������        ����                (           	      �       f        ��        ���� � �������������          ����                ,              >  |       f       ��        ���� � �������������          ����                0              \  �       f       ��        ���� � �������������          ����   	 
            4              z  �       f       ��       ���� � �������������          ����                8              �  0       f       ��       ���� � �������������          ����                <              �  l       f       ��       ���� � �������������          ����                @              �  �       f       ��       ���� � �������������          ����                D              �  �       f       ��       ���� � �������������          ����                H                        f       ��       ���� � �������������          ����                L              .  \       f	       ��       ���� � �������������          ����               '              �   �        4        ��        ���� � �������������          ����               +              �   �       4       ��        ���� � �������������          ����               /                       4       ��        ���� � �������������          ����  	 
            3              "  D       4       ��       ���� � �������������          ����               7              @  �       4       ��       ���� � �������������          ����               ;              ^  �       4       ��       ���� � �������������          ����               ?              |  �       4       ��       ���� � �������������          ����               C              �  4       4       ��       ���� � �������������          ����               G              �  p       4       ��       ���� � �������������          ����               K           	   �  �       4	       ��       ���� � �������������          ����                             ,  h       �        ��        ���� � �������������          ����               "              J  �       �       ��        ���� � �������������          ����               &              h  �       �       ��        ���� � �������������          ����  	 
            *              �         �       ��       ���� � �������������          ����               .              �  H       �       ��       ���� � �������������          ����               2           	   �  �       �       ��       ���� � �������������          ����               6           	   �  �       �       ��       ���� � �������������          ����               :           
   �  �       �       ��       ���� � �������������          ����               >           
     8       �       ��       ���� � �������������          ����               B              :  t       �	       ��       ���� � �������������          ����                          !   �  /       �        ��        ���� � �������������          ����                          (   �  �       �       ��        ���� � �������������          ����               #           )            �       ��        ���� � �������������          ����  	 
            '           )   *  T       �       ��       ���� � �������������          ����               +           *   H  �       �       ��       ���� � �������������          ����               /           +   f  �       �       ��       ���� � �������������          ����               3           +   �         �       ��       ���� � �������������          ����               7           ,   �  D       �       ��       ���� � �������������          ����               ;           ,   �  �       �       ��       ���� � �������������          ����               ?           -   �  �       �	       ��       ���� � �������������          ����                             �  F       f        ��        ���� � �������������          ����               #              �  �	       f       ��        ���� � �������������          ����   	            '              �  �	       f       ��        ���� � �������������          ����  
             +              
  
       f       ��       ���� � �������������          ����               /              (  P
       f       ��       ���� � �������������          ����               3              F  �
       f       ��       ���� � �������������          ����               7              d  �
       f       ��       ���� � �������������          ����               ;              �         f       ��       ���� � �������������          ����               ?              �  @       f       ��       ���� � �������������          ����               C              �  |       f	       ��       ���� � �������������          ����               2              @  �                 ��        ���� � �������������          ����               6               ^  �                ��        ���� � �������������          ����  	 
            :           !   |  �                ��        ���� � �������������          ����               >           !   �  4                ��       ���� � �������������          ����               B           "   �  p                ��       ���� � �������������          ����               F           #   �  �                ��       ���� � �������������          ����               J           #   �  �                ��       ���� � �������������          ����               N           $     $                ��       ���� � �������������          ����               R           $   0  `                ��       ���� � �������������          ����               V           %   N  �        	        ��       ���� � �������������          ����                /           �����  X       �      ��  ��        ���� � �������������          ����                3           ����  $       �     ��  ��        ���� � �������������          ����  	 
             7           ����0  `       �     ��  ��        ���� � �������������          ����                ;           ����N  �       �     ��  ��       ���� � �������������          ����                ?           ����l  �       �     ��  ��       ���� � �������������          ����                C           �����         �     ��  ��       ���� � �������������          ����                G           �����  P       �     ��  ��       ���� � �������������          ����                K           �����  �       �     ��  ��       ���� � �������������          ����                O           �����  �       �     ��  ��       ���� � �������������          ����                S           ����         �	     ��  ��       ���� � �������������          ����
                '           �����  t1       s      ��  ��        ���� � �������������          ����
                +           �����  <       s     ��  ��        ���� � �������������          ����
   	             /           �����  x       s     ��  ��        ���� � �������������          ����
  
              3           �����  �       s     ��  ��       ���� � �������������          ����
                7           �����  �       s     ��  ��       ���� � �������������          ����
                ;           ����  ,       s     ��  ��       ���� � �������������          ����
                ?           ����4  h       s     ��  ��       ���� � �������������          ����
                C           ����R  �       s     ��  ��       ���� � �������������          ����
                G           ����p  �       s     ��  ��       ���� � �������������          ����
                K           �����         s	     ��  ��       ���� � �������������            ��                3          �����
  �         �       �             ���� � �������������            ��                7          ����          �      �             ���� � �������������            ��   	             ;          ����,  X        �      �             ���� � �������������            ��  
              ?          ����J  �        �      �             ���� � �������������            ��                C          ����h  �        �      �             ���� � �������������            ��                G          �����          �      �             ���� � �������������            ��                K          �����  H        �      �             ���� � �������������            ��                O          �����  �        �      �             ���� � �������������            ��                S          �����  �        �      �             ���� � �������������            ��                W          �����  �        � 	     �             ���� � �������������          ����                9           ����0  �        �      ��  ��        ���� � �������������          ����                =           ����N  �"       �     ��  ��        ���� � �������������          ����  	 
             A           ����l  �"       �     ��  ��        ���� � �������������          ����                E           �����  #       �     ��  ��       ���� � �������������          ����                I           �����  P#       �     ��  ��       ���� � �������������          ����                M           �����  �#       �     ��  ��       ���� � �������������          ����                Q           �����  �#       �     ��  ��       ���� � �������������          ����                U           ����  $       �     ��  ��       ���� � �������������          ����                Y           ����   @$       �     ��  ��       ���� � �������������          ����                ]           ����>  |$       �	     ��  ��       ���� � �������������          ����	                           ����  .J             ��  ��        ���� � �������������          ����	                #           ����.  \            ��  ��        ���� � �������������          ����	                '           ����L  �            ��  ��        ���� � �������������          ����	  	 
             +           ����j  �            ��  ��       ���� � �������������          ����	                /           �����              ��  ��       ���� � �������������          ����	                3           �����  L            ��  ��       ���� � �������������          ����	                7           �����  �            ��  ��       ���� � �������������          ����	                ;           �����  �            ��  ��       ���� � �������������          ����	                ?           ����                ��  ��       ���� � �������������          ����	                C           ����  <       	     ��  ��       ���� � �������������          ����                7           �����  �        '      ��  ��        ���� � �������������          ����                ;           �����  |       '     ��  ��        ���� � �������������          ����  	 
             ?           �����  �       '     ��  ��        ���� � �������������          ����                C           �����  �       '     ��  ��       ���� � �������������          ����                G           ����  0        '     ��  ��       ���� � �������������          ����                K           ����6  l        '     ��  ��       ���� � �������������          ����                O           ����T  �        '     ��  ��       ���� � �������������          ����                S           ����r  �        '     ��  ��       ���� � �������������          ����                W           �����   !       '     ��  ��       ���� � �������������          ����                [           �����  \!       '	     ��  ��       ���� � �������������            g                             �����   �        #      ��( ��        ����   ����������������        ] g                           ����B  �        $      ��( ��        ����   ����������������        ^ g                          ����[  l        %      ��( ��        ����   ����������������        _ g                 &         ����'  �#        &      ��( ��         ����   ����������������        ` g                % .         �����
  �?        '      ��( ��!        ����   ����������������        a g                6 A + "       �����  �g        (      ��( ��"        ����   ����������������        b g                @ L 2 )       �����  �        )      ��( ��#        ����   ����������������        c g                W e = 1       ����U  ��        *      ��( ��$        ����   ����������������        d g                d s X :       �����  @<       +      ��( ��%        ����	   ����������������        e g                2*      �����  p�       ,      ��( ��&        ����
   ����������������        f g                � � � L       ����O.  �+       -      ��( ��'        ����   ����������������        g g                � � � U       �����6  �       .      ��( ��(        ����   ����������������        h g                ��(�       �����  <d
       /      ��( ��)        ����   ����������������        i g                � � � m       �����I  �O       0      ��( ��*        ����   ����������������        j g                � �       ����T  A       1      ��( ��+        ����   ����������������        k g                '<� �       ����A_  QS       2      ��( ��,        ����   ����������������        l g                K`� �       ����$k  ��       3      ��( ��-        ����   ����������������        m g                q��       �����w  ��       4      ��( ��.        ����   ����������������        n g                � � � b       �����?  }       5      ��( ��/        ����   ����������������        o g                ��D�       ������  �       6      ��( ��0        ����   ����������������        p g                �a      ������  ��       7      ��( ��1        ����   ����������������        q g                � � f A       �����&  ʨ       8      ��( ��2        ����   ����������������        r g                Mb�G      ����%�  x       9      ��( ��3        ����   ����������������        ����              $ 9           #   �  �       g        ��4        ���� � �������������          ����   	 
          ( =           %   �  �       g       ��4        ���� � �������������          ����              , A           '     Z       g       ��4        ���� � �������������          ����              0 E           )   Z         g       ��4       ���� � �������������          ����              4 I           *   �  �       g       ��4       ���� � �������������          ����              8 M           ,   �  v       g       ��4       ���� � �������������          ����              < Q           .     *       g       ��4       ���� � �������������          ����              @ U           0   J  �       g       ��4       ���� � �������������          ����              D Y           2   �  �       g       ��4       ���� � �������������          ����              H ]           3   �  F       g	       ��4       ���� � �������������          ����             $ 8              N  �       5        ��5        ���� � �������������          ����  	 
          ( <              �  �       5       ��5        ���� � �������������          ����             , @              �  R       5       ��5        ���� � �������������          ����             0 D                	       5       ��5       ���� � �������������          ����             4 H              >  �	       5       ��5       ���� � �������������          ����             8 L              z  n
       5       ��5       ���� � �������������          ����             < P              �  "       5       ��5       ���� � �������������          ����             @ T              �  �       5       ��5       ���� � �������������          ����             D X               .  �       5       ��5       ���� � �������������          ����             H \           !   j  >       5	       ��5       ���� � �������������          ����             $ /              �         �        ��6        ���� � �������������          ����  	 
          ( 3              �  �       �       ��6        ���� � �������������          ����             , 7              *  ~	       �       ��6        ���� � �������������          ����             0 ;              f  2
       �       ��6       ���� � �������������          ����             4 ?              �  �
       �       ��6       ���� � �������������          ����             8 C              �  �       �       ��6       ���� � �������������          ����             < G                N       �       ��6       ���� � �������������          ����             @ K           !   V         �       ��6       ���� � �������������          ����             D O           #   �  �       �       ��6       ���� � �������������          ����             H S           $   �  j       �	       ��6       ���� � �������������          ����             $ ,           G   V	         �        ��7        ���� � �������������          ����  	 
          ( 0           I   �	  �       �       ��7        ���� � �������������          ����             , 4           K   �	  j       �       ��7        ���� � �������������          ����             0 8           M   

         �       ��7       ���� � �������������          ����             4 <           N   F
  �       �       ��7       ���� � �������������          ����             8 @           P   �
  �       �       ��7       ���� � �������������          ����             < D           R   �
  :        �       ��7       ���� � �������������          ����             @ H           T   �
  �        �       ��7       ���� � �������������          ����             D L           V   6  �!       �       ��7       ���� � �������������          ����             H P           W   r  V"       �	       ��7       ���� � �������������          ����   	          $ 0           /   6  �       g        ��8        ���� � �������������          ����  
           ( 4           1   r  V       g       ��8        ���� � �������������          ����             , 8           3   �  
       g       ��8        ���� � �������������          ����             0 <           5   �  �       g       ��8       ���� � �������������          ����             4 @           6   &  r       g       ��8       ���� � �������������          ����             8 D           8   b  &       g       ��8       ���� � �������������          ����             < H           :   �  �       g       ��8       ���� � �������������          ����             @ L           <   �  �       g       ��8       ���� � �������������          ����             D P           >     B       g       ��8       ���� � �������������          ����             H T           ?   R  �       g	       ��8       ���� � �������������          ����  	 
          $ C           ;   �  R               ��9        ���� � �������������          ����             ( G           =                   ��9        ���� � �������������          ����             , K           ?   >  �              ��9        ���� � �������������          ����             0 O           A   z  n              ��9       ���� � �������������          ����             4 S           B   �  "              ��9       ���� � �������������          ����             8 W           D   �  �              ��9       ���� � �������������          ����             < [           F   .	  �              ��9       ���� � �������������          ����             @ _           H   j	  >              ��9       ���� � �������������          ����             D c           J   �	  �              ��9       ���� � �������������          ����             H g           K   �	  �       	       ��9       ���� � �������������          ����  	 
           $ @           ����z  n
       �      ��  ��:        ���� � �������������          ����              ( D           �����  "       �     ��  ��:        ���� � �������������          ����              , H           �����  �       �     ��  ��:        ���� � �������������          ����              0 L           ����.  �       �     ��  ��:       ���� � �������������          ����              4 P           ����j  >       �     ��  ��:       ���� � �������������          ����              8 T           �����  �       �     ��  ��:       ���� � �������������          ����              < X           �����  �       �     ��  ��:       ���� � �������������          ����              @ \           ����  Z       �     ��  ��:       ���� � �������������          ����              D `           ����Z         �     ��  ��:       ���� � �������������          ����              H d           �����  �       �	     ��  ��:       ���� � �������������          ����
   	           $ 8           ����  *       t      ��  ��;        ���� � �������������          ����
  
            ( <           ����B  �*       t     ��  ��;        ���� � �������������          ����
              , @           ����~  z+       t     ��  ��;        ���� � �������������          ����
              0 D           �����  .,       t     ��  ��;       ���� � �������������          ����
              4 H           �����  �,       t     ��  ��;       ���� � �������������          ����
              8 L           ����2  �-       t     ��  ��;       ���� � �������������          ����
              < P           ����n  J.       t     ��  ��;       ���� � �������������          ����
              @ T           �����  �.       t     ��  ��;       ���� � �������������          ����
              D X           �����  �/       t     ��  ��;       ���� � �������������          ����
              H \           ����"  f0       t	     ��  ��;       ���� � �������������           ��   	           $ D     (     ����v  b%        �       �     <        ���� � �������������           ��  
            ( H     (     �����  &        �      �     <        ���� � �������������           ��              , L     (     �����  �&        �      �     <        ���� � �������������           ��              0 P     (     ����*  ~'        �      �     <        ���� � �������������           ��              4 T     (     ����f  2(        �      �     <        ���� � �������������           ��              8 X     (     �����  �(        �      �     <        ���� � �������������           ��              < \     (     �����  �)        �      �     <        ���� � �������������           ��              @ `     (     ����  N*        �      �     <        ���� � �������������           ��              D d     (     ����V  +        �      �     <        ���� � �������������           ��              H h     (     �����  �+        � 	     �     <        ���� � �������������          ����  	 
           $ J           �����  "8       �      ��  ��=        ���� � �������������          ����              ( N           �����  �8       �     ��  ��=        ���� � �������������          ����              , R           ����.  �9       �     ��  ��=        ���� � �������������          ����              0 V           ����j  >:       �     ��  ��=       ���� � �������������          ����              4 Z           �����  �:       �     ��  ��=       ���� � �������������          ����              8 ^           �����  �;       �     ��  ��=       ���� � �������������          ����              < b           ����  Z<       �     ��  ��=       ���� � �������������          ����              @ f           ����Z  =       �     ��  ��=       ���� � �������������          ����              D j           �����  �=       �     ��  ��=       ���� � �������������          ����              H n           �����  v>       �	     ��  ��=       ���� � �������������          ����	              $ 0           �����  �.             ��  ��>        ���� � �������������          ����	  	 
           ( 4           �����  v/            ��  ��>        ���� � �������������          ����	              , 8           ����  *0            ��  ��>        ���� � �������������          ����	              0 <           ����J  �0            ��  ��>       ���� � �������������          ����	              4 @           �����  �1            ��  ��>       ���� � �������������          ����	              8 D           �����  F2            ��  ��>       ���� � �������������          ����	              < H           �����  �2            ��  ��>       ���� � �������������          ����	              @ L           ����:  �3            ��  ��>       ���� � �������������          ����	              D P           ����v  b4            ��  ��>       ���� � �������������          ����	              H T           �����  5       	     ��  ��>       ���� � �������������          ����  	 
           $ H           ����&  r3       (      ��  ��?        ���� � �������������          ����              ( L           ����b  &4       (     ��  ��?        ���� � �������������          ����              , P           �����  �4       (     ��  ��?        ���� � �������������          ����              0 T           �����  �5       (     ��  ��?       ���� � �������������          ����              4 X           ����  B6       (     ��  ��?       ���� � �������������          ����              8 \           ����R  �6       (     ��  ��?       ���� � �������������          ����              < `           �����  �7       (     ��  ��?       ���� � �������������          ����              @ d           �����  ^8       (     ��  ��?       ���� � �������������          ����              D h           ����  9       (     ��  ��?       ���� � �������������          ����              H l           ����B  �9       (	     ��  ��?       ���� � �������������          ����              5 I          N   �  �       h        ��@        ���� � ������������          ����              : N !         R     0        h       ��@        ���� � ������������          ����              ? S $         V   f  �!       h       ��@        ���� � ������������          ����              D X '         Y   �   #       h       ��@       ���� � ������������          ����              I ] *         ]   	  h$       h       ��@       ���� � ������������          ����              N b -         `   t	  �%       h       ��@       ���� � ������������          ����              S g 0         d   �	  8'       h       ��@       ���� � ������������          ����              X l 3         h   (
  �(       h       ��@       ���� � ������������          ����              ] q 6         k   �
  *       h       ��@       ���� � ������������          ����              b v 9         o   �
  p+       h	       ��@       ���� � ������������          ����             5 H          6   Z  h       6        ��A        ���� � ������������         ����             : M !         :   �  �       6       ��A        ���� � ������������         ����             ? R $         >     8       6       ��A        ���� � ������������         ����             D W '         A   h  �       6       ��A       ���� � ������������         ����             I \ *         E   �         6       ��A       ���� � ������������         ����             N a -         H     p       6       ��A       ���� � ������������         ����             S f 0         L   v  �       6       ��A       ���� � ������������         ����             X k 3         P   �  @       6       ��A       ���� � ������������         ����             ] p 6         S   *  �        6       ��A       ���� � ������������         ����             b u 9         W   �  "       6	       ��A       ���� � ������������          ����             5 ?          :   �  �       �        ��B        ���� � ������������         ����             : D !         >     `       �       ��B        ���� � ������������         ����             ? I $         B   r  �       �       ��B        ���� � ������������         ����             D N '         E   �  0       �       ��B       ���� � ������������         ����             I S *         I   &  �       �       ��B       ���� � ������������         ����             N X -         L   �          �       ��B       ���� � ������������         ����             S ] 0         P   �  h       �       ��B       ���� � ������������         ����             X b 3         T   4  �        �       ��B       ���� � ������������         ����             ] g 6         W   �  8"       �       ��B       ���� � ������������         ����             b l 9         [   �  �#       �	       ��B       ���� � ������������          ����             5 <          ~   b  �1       �        ��C        ���� � ������������         ����             : A !         �   �  �2       �       ��C        ���� � ������������         ����             ? F $         �     X4       �       ��C        ���� � ������������         ����             D K '         �   p  �5       �       ��C       ���� � ������������         ����             I P *         �   �  (7       �       ��C       ���� � ������������         ����             N U -         �   $  �8       �       ��C       ���� � ������������         ����             S Z 0         �   ~  �9       �       ��C       ���� � ������������         ����             X _ 3         �   �  `;       �       ��C       ���� � ������������         ����             ] d 6         �   2  �<       �       ��C       ���� � ������������         ����             b i 9         �   �  0>       �	       ��C       ���� � ������������          ����             5 @          ^   B	  %       h        ��D        ���� � ������������         ����             : E !         b   �	  p&       h       ��D        ���� � ������������         ����             ? J $         f   �	  �'       h       ��D        ���� � ������������         ����             D O '         i   P
  @)       h       ��D       ���� � ������������         ����             I T *         m   �
  �*       h       ��D       ���� � ������������         ����             N Y -         p     ,       h       ��D       ���� � ������������         ����             S ^ 0         t   ^  x-       h       ��D       ���� � ������������         ����             X c 3         x   �  �.       h       ��D       ���� � ������������         ����             ] h 6         {     H0       h       ��D       ���� � ������������         ����              b m 9            l  �1       h	       ��D       ���� � ������������         ����             5 S          n   �
  H+               ��E        ���� � ������������         ����             : X !         r   ,  �,              ��E        ���� � ������������         ����             ? ] $         v   �  .              ��E        ���� � ������������         ����             D b '         y   �  �/              ��E       ���� � ������������         ����             I g *         }   :  �0              ��E       ���� � ������������         ����             N l -         �   �  P2              ��E       ���� � ������������         ����             S q 0         �   �  �3              ��E       ���� � ������������         ����             X v 3         �   H   5              ��E       ���� � ������������         ����             ] { 6         �   �  �6              ��E       ���� � ������������         ����    !          b � 9         �   �  �7       	       ��E       ���� � ������������         ����              5 P          �����         �      ��  ��F        ���� � ������������         ����              : U !         �����  �       �     ��  ��F        ���� � ������������         ����              ? Z $         ����:  �       �     ��  ��F        ���� � ������������         ����              D _ '         �����  P       �     ��  ��F       ���� � ������������         ����              I d *         �����  �       �     ��  ��F       ���� � ������������         ����              N i -         ����H   !       �     ��  ��F       ���� � ������������         ����              S n 0         �����  �"       �     ��  ��F       ���� � ������������         ����              X s 3         �����  �#       �     ��  ��F       ���� � ������������         ����              ] x 6         ����V	  X%       �     ��  ��F       ���� � ������������         ����    !           b } 9         �����	  �&       �	     ��  ��F       ���� � ������������         ����
              5 H          ����  HD       u      ��  ��G        ���� � ������������         ����
              : M !         ����l  �E       u     ��  ��G        ���� � ������������         ����
              ? R $         �����  G       u     ��  ��G        ���� � ������������         ����
              D W '         ����   �H       u     ��  ��G       ���� � ������������         ����
              I \ *         ����z  �I       u     ��  ��G       ���� � ������������         ����
              N a -         �����  PK       u     ��  ��G       ���� � ������������         ����
              S f 0         ����.  �L       u     ��  ��G       ���� � ������������         ����
              X k 3         �����   N       u     ��  ��G       ���� � ������������         ����
              ] p 6         �����  �O       u     ��  ��G       ���� � ������������         ����
               b u 9         ����<  �P       u	     ��  ��G       ���� � ������������          ��              5 T    2     �����  >        �       �     H        ���� � ������������          ��              : Y !   2     �����  p?        �      �     H        ���� � ������������          ��              ? ^ $   2     ����6  �@        �      �     H        ���� � ������������          ��              D c '   2     �����  @B        �      �     H        ���� � ������������          ��              I h *   2     �����  �C        �      �     H        ���� � ������������          ��              N m -   2     ����D  E        �      �     H        ���� � ������������          ��              S r 0   2     �����  xF        �      �     H        ���� � ������������          ��              X w 3   2     �����  �G        �      �     H        ���� � ������������          ��              ] | 6   2     ����R  HI        �      �     H        ���� � ������������          ��               b � 9   2     �����  �J        � 	     �     H        ���� � ������������         ����              5 Z          �����  W       �      ��  ��I        ���� � ������������	         ����              : _ !         ����  pX       �     ��  ��I        ���� � ������������	         ����              ? d $         ����v  �Y       �     ��  ��I        ���� � ������������	         ����              D i '         �����  @[       �     ��  ��I       ���� � ������������	         ����              I n *         ����*  �\       �     ��  ��I       ���� � ������������	         ����              N s -         �����  ^       �     ��  ��I       ���� � ������������	         ����              S x 0         �����  x_       �     ��  ��I       ���� � ������������	         ����              X } 3         ����8  �`       �     ��  ��I       ���� � ������������	         ����              ] � 6         �����  Hb       �     ��  ��I       ���� � ������������	         ����    !           b � 9         �����  �c       �	     ��  ��I       ���� � ������������	         ����	              5 @          �����  �J             ��  ��J        ���� � ������������
         ����	              : E !         �����  �K            ��  ��J        ���� � ������������
         ����	              ? J $         ����V  XM            ��  ��J        ���� � ������������
         ����	              D O '         �����  �N            ��  ��J       ���� � ������������
         ����	              I T *         ����
  (P            ��  ��J       ���� � ������������
         ����	              N Y -         ����d  �Q            ��  ��J       ���� � ������������
         ����	              S ^ 0         �����  �R            ��  ��J       ���� � ������������
         ����	              X c 3         ����  `T            ��  ��J       ���� � ������������
         ����	              ] h 6         ����r  �U            ��  ��J       ���� � ������������
         ����	              b m 9         �����  0W       	     ��  ��J       ���� � ������������
         ����              5 X          ����2  �P       )      ��  ��K        ���� � ������������         ����              : ] !         �����  0R       )     ��  ��K        ���� � ������������         ����              ? b $         �����  �S       )     ��  ��K        ���� � ������������         ����              D g '         ����@   U       )     ��  ��K       ���� � ������������         ����              I l *         �����  hV       )     ��  ��K       ���� � ������������         ����              N q -         �����  �W       )     ��  ��K       ���� � ������������         ����              S v 0         ����N  8Y       )     ��  ��K       ���� � ������������         ����              X { 3         �����  �Z       )     ��  ��K       ���� � ������������         ����              ] � 6         ����  \       )     ��  ��K       ���� � ������������         ����    !           b � 9         ����\  p]       )	     ��  ��K       ���� � ������������          ����              O b &        �   D  T=       i        ��L        ���� � ������������         ����              T g )        �   �  �?       i       ��L        ���� � ������������         ����              Y l ,         �   4  B       i       ��L        ���� � ������������         ����              ^ q / #       �   �  \D       i       ��L       ���� � ������������         ����              c v 2 &       �   $  �F       i       ��L       ���� � ������������         ����              h { 5 )       �   �  I       i       ��L       ���� � ������������         ����              m � 8 ,       �     dK       i       ��L       ���� � ������������         ����              r � ; /       �   �  �M       i       ��L       ���� � ������������         ����     !          w � > 2       �     P       i       ��L       ���� � ������������         ����   " #          | � A 5       �   |  lR       i	       ��L       ���� � ������������         ����             O a &           �	  �1       7        ��M        ���� � ������������         ����             T f )        �   d
  �3       7       ��M        ���� � ������������         ����             Y k ,         �   �
  L6       7       ��M        ���� � ������������         ����             ^ p / #       �   T  �8       7       ��M       ���� � ������������         ����             c u 2 &       �   �  �:       7       ��M       ���� � ������������         ����             h z 5 )       �   D  T=       7       ��M       ���� � ������������         ����             m  8 ,       �   �  �?       7       ��M       ���� � ������������         ����             r � ; /       �   4  B       7       ��M       ���� � ������������         ����    !          w � > 2       �   �  \D       7       ��M       ���� � ������������         ����  " #          | � A 5       �   $  �F       7	       ��M       ���� � ������������          ����             O X &        �   P
  �3       �        ��N        ���� � ������������         ����             T ] )        �   �
  �5       �       ��N        ���� � ������������         ����             Y b ,         �   @  @8       �       ��N        ���� � ������������         ����             ^ g / #       �   �  �:       �       ��N       ���� � ������������         ����             c l 2 &       �   0  �<       �       ��N       ���� � ������������         ����             h q 5 )       �   �  H?       �       ��N       ���� � ������������         ����             m v 8 ,       �      �A       �       ��N       ���� � ������������         ����             r { ; /       �   �  �C       �       ��N       ���� � ������������         ����    !          w � > 2       �     PF       �       ��N       ���� � ������������         ����  " #          | � A 5       �   �  �H       �	       ��N       ���� � ������������          ����             O U &        �   �  �T       �        ��O        ���� � ������������         ����             T Z )        �   l  W       �       ��O        ���� � ������������         ����             Y _ ,         �   �  tY       �       ��O        ���� � ������������         ����             ^ d / #       �   \  �[       �       ��O       ���� � ������������         ����             c i 2 &       �   �  $^       �       ��O       ���� � ������������         ����             h n 5 )       �   L  |`       �       ��O       ���� � ������������         ����             m s 8 ,       �   �  �b       �       ��O       ���� � ������������         ����             r x ; /         <  ,e       �       ��O       ���� � ������������         ����    !          w } > 2       	  �  �g       �       ��O       ���� � ������������         ����  " #          | � A 5         ,  �i       �	       ��O       ���� � ������������          ����             O Y &        �   �  $E       i        ��P        ���� � ������������         ����             T ^ )        �   L  |G       i       ��P        ���� � ������������         ����             Y c ,         �   �  �I       i       ��P        ���� � ������������         ����             ^ h / #       �   <  ,L       i       ��P       ���� � ������������         ����             c m 2 &       �   �  �N       i       ��P       ���� � ������������         ����             h r 5 )       �   ,  �P       i       ��P       ���� � ������������         ����             m w 8 ,       �   �  4S       i       ��P       ���� � ������������         ����              r | ; /       �     �U       i       ��P       ���� � ������������         ����  ! "          w � > 2       �   �  �W       i       ��P       ���� � ������������         ����  # $          | � A 5       �     <Z       i	       ��P       ���� � ������������         ����             O l &        �   d  �L               ��Q        ���� � ������������         ����             T q )        �   �  LO              ��Q        ���� � ������������         ����             Y v ,         �   T  �Q              ��Q        ���� � ������������         ����             ^ { / #       �   �  �S              ��Q       ���� � ������������         ����             c � 2 &       �   D  TV              ��Q       ���� � ������������         ����             h � 5 )       �   �  �X              ��Q       ���� � ������������         ����             m � 8 ,       �   4  [              ��Q       ���� � ������������         ����    !          r � ; /       �   �  \]              ��Q       ���� � ������������         ����  " #          w � > 2       �   $  �_              ��Q       ���� � ������������         ����  $ %          | � A 5       �   �  b       	       ��Q       ���� � ������������         ����              O i &        ����  x7       �      ��  ��R        ���� � ������������         ����              T n )        �����  �9       �     ��  ��R        ���� � ������������         ����              Y s ,         ����  (<       �     ��  ��R        ���� � ������������         ����              ^ x / #       �����  �>       �     ��  ��R       ���� � ������������         ����              c } 2 &       �����  �@       �     ��  ��R       ���� � ������������         ����              h � 5 )       ����p  0C       �     ��  ��R       ���� � ������������         ����              m � 8 ,       �����  �E       �     ��  ��R       ���� � ������������         ����    !           r � ; /       ����`  �G       �     ��  ��R       ���� � ������������         ����  " #           w � > 2       �����  8J       �     ��  ��R       ���� � ������������         ����  $ %           | � A 5       ����P  �L       �	     ��  ��R       ���� � ������������         ����
              O a &        �����  4l       v      ��  ��S        ���� � ������������         ����
              T f )        ����  �n       v     ��  ��S        ���� � ������������         ����
              Y k ,         �����  �p       v     ��  ��S        ���� � ������������         ����
              ^ p / #       ����  <s       v     ��  ��S       ���� � ������������         ����
              c u 2 &       �����  �u       v     ��  ��S       ���� � ������������         ����
              h z 5 )       �����  �w       v     ��  ��S       ���� � ������������         ����
              m  8 ,       ����t  Dz       v     ��  ��S       ���� � ������������         ����
               r � ; /       �����  �|       v     ��  ��S       ���� � ������������         ����
  ! "           w � > 2       ����d  �~       v     ��  ��S       ���� � ������������         ����
  # $           | � A 5       �����  L�       v	     ��  ��S       ���� � ������������         	 ��              O m &  <     ����  dd        �       �     T        ���� � ������������         	 ��              T r )  <     �����  �f        �      �     T        ���� � ������������         	 ��              Y w ,   <     ����  i        �      �     T        ���� � ������������         	 ��              ^ | / # <     ����|  lk        �      �     T        ���� � ������������         	 ��              c � 2 & <     �����  �m        �      �     T        ���� � ������������         	 ��              h � 5 ) <     ����l  p        �      �     T        ���� � ������������         	 ��              m � 8 , <     �����  tr        �      �     T        ���� � ������������         	 ��               r � ; / <     ����\  �t        �      �     T        ���� � ������������         	 ��  ! "           w � > 2 <     �����  $w        �      �     T        ���� � ������������         	 ��  # $           | � A 5 <     ����L  |y        � 	     �     T        ���� � ������������         ����              O s &        ����T  ��       �      ��  ��U        ���� � ������������         ����              T x )        �����  ��       �     ��  ��U        ���� � ������������         ����              Y } ,         ����D  T�       �     ��  ��U        ���� � ������������         ����              ^ � / #       �����  ��       �     ��  ��U       ���� � ������������         ����              c � 2 &       ����4  �       �     ��  ��U       ���� � ������������         ����              h � 5 )       �����  \�       �     ��  ��U       ���� � ������������         ����              m � 8 ,       ����$  ��       �     ��  ��U       ���� � ������������         ����    !           r � ; /       �����  �       �     ��  ��U       ���� � ������������         ����  " #           w � > 2       ����  d�       �     ��  ��U       ���� � ������������         ����  $ %           | � A 5       �����  ��       �	     ��  ��U       ���� � ������������         ����	              O Y &        ����4  t             ��  ��V        ���� � ������������         ����	              T ^ )        �����  \v            ��  ��V        ���� � ������������         ����	              Y c ,         ����$  �x            ��  ��V        ���� � ������������         ����	              ^ h / #       �����  {            ��  ��V       ���� � ������������         ����	              c m 2 &       ����  d}            ��  ��V       ���� � ������������         ����	              h r 5 )       �����  �            ��  ��V       ���� � ������������         ����	              m w 8 ,       ����  �            ��  ��V       ���� � ������������         ����	              r | ; /       ����|  l�            ��  ��V       ���� � ������������         ����	    !           w � > 2       �����  Ć            ��  ��V       ���� � ������������         ����	  " #           | � A 5       ����l  �       	     ��  ��V       ���� � ������������         ����              O q &        �����  �{       *      ��  ��W        ���� � ������������         ����              T v )        ����<  ,~       *     ��  ��W        ���� � ������������         ����              Y { ,         �����  ��       *     ��  ��W        ���� � ������������         ����              ^ � / #       ����,  ܂       *     ��  ��W       ���� � ������������         ����              c � 2 &       �����  4�       *     ��  ��W       ���� � ������������         ����              h � 5 )       ����  ��       *     ��  ��W       ���� � ������������         ����              m � 8 ,       �����  �       *     ��  ��W       ���� � ������������         ����    !           r � ; /       ����  <�       *     ��  ��W       ���� � ������������         ����  " #           w � > 2       �����  ��       *     ��  ��W       ���� � ������������         ����  $ %           | � A 5       �����  �       *	     ��  ��W       ���� � ������������          ����              h z - !         \  (n       j        ��X        ���� � ������������         ����              m  0 $       #  �  �q       j       ��X        ���� � ������������         ����              r � 3 '       ,  �  0u       j       ��X        ���� � ������������         ����              w � 6 *       5    �x       j       ��X       ���� � ������������         ����              | � 9 -       >  �  8|       j       ��X       ���� � ������������         ����              � � < 0       G  J  �       j       ��X       ���� � ������������         ����     !          � � ? 3       P  �  @�       j       ��X       ���� � ������������         ����   " #          � � B 6       Y  v  Ć       j       ��X       ���� � ������������         ����   $ %          � � E 9       b    H�    
   j       ��X       ���� � ������������         ����   & '          � � H <       k  �  ̍    	   j	       ��X       ���� � ������������         ����             h y - !       �     `       8        ��Y        ���� � ������������         ����             m ~ 0 $       �   �  �c       8       ��Y        ���� � ������������         ����             r � 3 '         0   g       8       ��Y        ���� � ������������         ����             w � 6 *         �  �j       8       ��Y       ���� � ������������         ����             | � 9 -         \  (n       8       ��Y       ���� � ������������         ����             � � < 0       #  �  �q       8       ��Y       ���� � ������������         ����    !          � � ? 3       ,  �  0u       8       ��Y       ���� � ������������         ����  " #          � � B 6       5    �x       8       ��Y       ���� � ������������         ����  $ %          � � E 9       >  �  8|    
   8       ��Y       ���� � ������������         ����  & '          � � H <       G  J  �    	   8	       ��Y       ���� � ������������          ����             h p - !       �   h  pb       �        ��Z        ���� � ������������         ����             m u 0 $         �  �e       �       ��Z        ���� � ������������         ����             r z 3 '         �  xi       �       ��Z        ���� � ������������         ����             w  6 *         *  �l       �       ��Z       ���� � ������������         ����             | � 9 -          �  �p       �       ��Z       ���� � ������������         ����             � � < 0       )  V  t       �       ��Z       ���� � ������������         ����    !          � � ? 3       2  �  �w       �       ��Z       ���� � ������������         ����  " #          � � B 6       ;  �  {       �       ��Z       ���� � ������������         ����  $ %          � � E 9       D    �~    
   �       ��Z       ���� � ������������         ����  & '          � � H <       M  �  �    	   �	       ��Z       ���� � ������������          ����             h m - !       b    H�       �        ��[        ���� � ������������         ����             m r 0 $       k  �  ̍       �       ��[        ���� � ������������         ����             r w 3 '       t  8  P�       �       ��[        ���� � ������������         ����             w | 6 *       }  �  Ԕ       �       ��[       ���� � ������������         ����             | � 9 -       �  d  X�       �       ��[       ���� � ������������         ����             � � < 0       �  �  ܛ       �       ��[       ���� � ������������         ����    !          � � ? 3       �  �  `�       �       ��[       ���� � ������������         ����  " #          � � B 6       �  &  �       �       ��[       ���� � ������������         ����  $ %          � � E 9       �  �  h�    
   �       ��[       ���� � ������������         ����  & '          � � H <       �  R  �    	   �	       ��[       ���� � ������������          ����             h q - !       2  �  �w       j        ��\        ���� � ������������         ����             m v 0 $       ;  �  {       j       ��\        ���� � ������������         ����             r { 3 '       D    �~       j       ��\        ���� � ������������         ����             w � 6 *       M  �  �       j       ��\       ���� � ������������         ����             | � 9 -       V  D  ��       j       ��\       ���� � ������������         ����              � � < 0       _  �  �       j       ��\       ���� � ������������         ����  ! "          � � ? 3       h  p  ��       j       ��\       ���� � ������������         ����  # $          � � B 6       q    $�       j       ��\       ���� � ������������         ����  % &          � � E 9       z  �  ��    
   j       ��\       ���� � ������������         ����  ' (          � � H <       �  2  ,�    	   j	       ��\       ���� � ������������         ����             h � - !       J  |  �               ��]        ���� � ������������         ����             m � 0 $       S    l�              ��]        ���� � ������������         ����             r � 3 '       \  �  ��              ��]        ���� � ������������         ����             w � 6 *       e  >  t�              ��]       ���� � ������������         ����             | � 9 -       n  �  ��              ��]       ���� � ������������         ����    !          � � < 0       w  j  |�              ��]       ���� � ������������         ����  " #          � � ? 3       �      �              ��]       ���� � ������������         ����  $ %          � � B 6       �  �  ��              ��]       ���� � ������������         ����  & '          � � E 9       �  ,  �    
          ��]       ���� � ������������         ����  ( )          � � H <       �  �  ��    	   	       ��]       ���� � ������������         ����              h � - !       ����0   g       �      ��  ��^        ���� � ������������         ����              m � 0 $       �����  �j       �     ��  ��^        ���� � ������������         ����              r � 3 '       ����\  (n       �     ��  ��^        ���� � ������������         ����              w � 6 *       �����  �q       �     ��  ��^       ���� � ������������         ����              | � 9 -       �����  0u       �     ��  ��^       ���� � ������������         ����    !           � � < 0       ����  �x       �     ��  ��^       ���� � ������������         ����  " #           � � ? 3       �����  8|       �     ��  ��^       ���� � ������������         ����  $ %           � � B 6       ����J  �       �     ��  ��^       ���� � ������������         ����  & '           � � E 9       �����  @�    
   �     ��  ��^       ���� � ������������         ����  ( )           � � H <       ����v  Ć    	   �	     ��  ��^       ���� � ������������         ����
              h y - !       �����  h�       w      ��  ��_        ���� � ������������         ����
              m ~ 0 $       ����R  �       w     ��  ��_        ���� � ������������         ����
              r � 3 '       �����  p�       w     ��  ��_        ���� � ������������         ����
              w � 6 *       ����~  ��       w     ��  ��_       ���� � ������������         ����
              | � 9 -       ����  x�       w     ��  ��_       ���� � ������������         ����
               � � < 0       �����  ��       w     ��  ��_       ���� � ������������         ����
  ! "           � � ? 3       ����@  ��       w     ��  ��_       ���� � ������������         ����
  # $           � � B 6       �����  �       w     ��  ��_       ���� � ������������         ����
  % &           � � E 9       ����l   ��    
   w     ��  ��_       ���� � ������������         ����
  ' (           � � H <       ����!  �    	   w	     ��  ��_       ���� � ������������         
 ��              h � - ! F     ����,  �        �       �     `        ���� � ������������          
 ��              m � 0 $ F     �����  ��        �      �     `        ���� � ������������          
 ��              r � 3 ' F     ����X  �        �      �     `        ���� � ������������           ��              w � 6 * F     �����  ��        �      �     `        ���� � ������������           ��              | � 9 - F     �����  �        �      �     `        ���� � ������������           ��               � � < 0 F     ����  ��        �      �     `        ���� � ������������           ��  ! "           � � ? 3 F     �����   �        �      �     `        ���� � ������������           ��  # $           � � B 6 F     ����F  ��        �      �     `        ���� � ������������           ��  % &           � � E 9 F     �����  (�        �      �     `        ���� � ������������           ��  ' (           � � H < F     ����r  ��        � 	     �     `        ���� � ������������          ����              h � - !       ����l   ��       �      ��  ��a        ���� � ������������!         ����              m � 0 $       ����!  �       �     ��  ��a        ���� � ������������!         ����              r � 3 '       �����!  ��       �     ��  ��a        ���� � ������������!         ����              w � 6 *       ����."  �       �     ��  ��a       ���� � ������������!         ����              | � 9 -       �����"  ��       �     ��  ��a       ���� � ������������!         ����    !           � � < 0       ����Z#  �       �     ��  ��a       ���� � ������������!         ����  " #           � � ? 3       �����#  ��       �     ��  ��a       ���� � ������������!         ����  $ %           � � B 6       �����$  $�       �     ��  ��a       ���� � ������������!         ����  & '           � � E 9       ����%  ��    
   �     ��  ��a       ���� � ������������!         ����  ( )           � � H <       �����%  ,�    	   �	     ��  ��a       ���� � ������������!         ����	              h q - !       ����L  ȯ             ��  ��b        ���� � ������������"         ����	              m v 0 $       �����  L�            ��  ��b        ���� � ������������"         ����	              r { 3 '       ����x  ж            ��  ��b        ���� � ������������"         ����	              w � 6 *       ����  T�            ��  ��b       ���� � ������������"         ����	              | � 9 -       �����  ؽ            ��  ��b       ���� � ������������"         ����	              � � < 0       ����:   \�            ��  ��b       ���� � ������������"         ����	    !           � � ? 3       �����   ��            ��  ��b       ���� � ������������"         ����	  " #           � � B 6       ����f!  d�            ��  ��b       ���� � ������������"         ����	  $ %           � � E 9       �����!  ��    
        ��  ��b       ���� � ������������"         ����	  & '           � � H <       �����"  l�    	   	     ��  ��b       ���� � ������������"         ����              h � - !       �����  (�       +      ��  ��c        ���� � ������������#         ����              m � 0 $       ����r  ��       +     ��  ��c        ���� � ������������#         ����              r � 3 '       ����   0�       +     ��  ��c        ���� � ������������#         ����              w � 6 *       �����   ��       +     ��  ��c       ���� � ������������#         ����              | � 9 -       ����4!  8�       +     ��  ��c       ���� � ������������#         ����    !           � � < 0       �����!  ��       +     ��  ��c       ���� � ������������#         ����  " #           � � ? 3       ����`"  @�       +     ��  ��c       ���� � ������������#         ����  $ %           � � B 6       �����"  ��       +     ��  ��c       ���� � ������������#         ����  & '           � � E 9       �����#  H�    
   +     ��  ��c       ���� � ������������#         ����  ( )           � � H <       ����"$  ��    	   +	     ��  ��c       ���� � ������������#          ����              � � 4 (       �  �  ֵ       k        ��d        ���� � ������������$         ����              � � 7 +       �  �  º       k       ��d        ���� � ������������$         ����              � � : .       �  b  ��       k       ��d        ���� � ������������$         ����              � � = 1       �    ��       k       ��d       ���� � ������������$         ����               � � @ 4         �  ��       k       ��d       ���� � ������������$         ����   " #          � � C 7         ~  r�       k       ��d       ���� � ������������$         ����   $ %          � � F :         2  ^�       k       ��d       ���� � ������������$         ����   & '          � � I =       )  �  J�    	   k       ��d       ���� � ������������$         ����   ( )          � � L @       6  �  6�       k       ��d       ���� � ������������$         ����   * +          � � O C       B  N   "�       k	       ��d       ���� � ������������$         ����             � � 4 (       �  �  n�       9        ��e        ���� � ������������%         ����             � � 7 +       �  V  Z�       9       ��e        ���� � ������������%         ����             � � : .       �  
  F�       9       ��e        ���� � ������������%         ����             � � = 1       �  �  2�       9       ��e       ���� � ������������%         ����              � � @ 4       �  r  �       9       ��e       ���� � ������������%         ����  " #          � � C 7       �  &  
�       9       ��e       ���� � ������������%         ����  $ %          � � F :       �  �  ��       9       ��e       ���� � ������������%         ����  & '          � � I =       �  �  ��    	   9       ��e       ���� � ������������%         ����  ( )          � � L @         B  ��       9       ��e       ���� � ������������%         ����  * +          � � O C         �  ��       9	       ��e       ���� � ������������%          ����             � � 4 (       �    *�       �        ��f        ���� � ������������&         ����             � � 7 +       �  �  �       �       ��f        ���� � ������������&         ����             � � : .       �  n  �       �       ��f        ���� � ������������&         ����             � � = 1       �  "  �       �       ��f       ���� � ������������&         ����              � � @ 4       �  �  ڻ       �       ��f       ���� � ������������&         ����  " #          � � C 7       �  �  ��       �       ��f       ���� � ������������&         ����  $ %          � � F :       �  >  ��       �       ��f       ���� � ������������&         ����  & '          � � I =         �  ��    	   �       ��f       ���� � ������������&         ����  ( )          � � L @         �  ��       �       ��f       ���� � ������������&         ����  * +          � � O C         Z  v�       �	       ��f       ���� � ������������&          ����             � � 4 (       %  �  ��       �        ��g        ���� � ������������'         ����             � � 7 +       2  ^  ��       �       ��g        ���� � ������������'         ����             � � : .       >     ~�       �       ��g        ���� � ������������'         ����             � � = 1       K  �   j�       �       ��g       ���� � ������������'         ����              � � @ 4       W  z!  V�       �       ��g       ���� � ������������'         ����  " #          � � C 7       d  ."  B�       �       ��g       ���� � ������������'         ����  $ %          � � F :       q  �"  .�       �       ��g       ���� � ������������'         ����  & '          � � I =       }  �#  �    	   �       ��g       ���� � ������������'         ����  ( )          � � L @       �  J$  �       �       ��g       ���� � ������������'         ����  * +          � � O C       �  �$  �      �	       ��g       ���� � ������������'          ����             � � 4 (       �  �  ��       k        ��h        ���� � ������������(         ����             � � 7 +       �  >  ��       k       ��h        ���� � ������������(         ����             � � : .         �  ��       k       ��h        ���� � ������������(         ����             � � = 1         �  ��       k       ��h       ���� � ������������(         ����    !          � � @ 4         Z  v�       k       ��h       ���� � ������������(         ����  # $          � � C 7       ,    b�       k       ��h       ���� � ������������(         ����  % &          � � F :       9  �  N�       k       ��h       ���� � ������������(         ����  ' (          � � I =       E  v   :�    	   k       ��h       ���� � ������������(         ����  ) *          � � L @       R  *!  &�       k       ��h       ���� � ������������(         ����  + ,          � � O C       ^  �!  �       k	       ��h       ���� � ������������(         ����             � � 4 (       	    ��               ��i        ���� � ������������)         ����             � � 7 +         �  ��              ��i        ���� � ������������)         ����             � � : .       "  �  ��              ��i        ���� � ������������)         ����              � � = 1       /  6  z�              ��i       ���� � ������������)         ����  ! "          � � @ 4       ;  �  f�              ��i       ���� � ������������)         ����  $ %          � � C 7       H  �   R�              ��i       ���� � ������������)         ����  & '          � � F :       U  R!  >�              ��i       ���� � ������������)         ����  ( )          � � I =       a  "  *�    	          ��i       ���� � ������������)         ����  * +          � � L @       n  �"  �              ��i       ���� � ������������)         ����  , -          � � O C       z  n#  �       	       ��i       ���� � ������������)         ����              � � 4 (       �����  ��       �      ��  ��j        ���� � ������������*         ����              � � 7 +       �����  ��       �     ��  ��j        ���� � ������������*         ����              � � : .       ����6  z�       �     ��  ��j        ���� � ������������*         ����               � � = 1       �����  f�       �     ��  ��j       ���� � ������������*         ����  ! "           � � @ 4       �����  R�       �     ��  ��j       ���� � ������������*         ����  $ %           � � C 7       ����R  >�       �     ��  ��j       ���� � ������������*         ����  & '           � � F :       ����  *�       �     ��  ��j       ���� � ������������*         ����  ( )           � � I =       �����  �    	   �     ��  ��j       ���� � ������������*         ����  * +           � � L @       ����n  �       �     ��  ��j       ���� � ������������*         ����  , -           � � O C       ����"  ��       �	     ��  ��j       ���� � ������������*         ����
              � � 4 (       ����Z#  v�       x      ��  ��k        ���� � ������������+         ����
              � � 7 +       ����$  b�       x     ��  ��k        ���� � ������������+         ����
              � � : .       �����$  N      x     ��  ��k        ���� � ������������+         ����
              � � = 1       ����v%  :      x     ��  ��k       ���� � ������������+         ����
    !           � � @ 4       ����*&  &      x     ��  ��k       ���� � ������������+         ����
  # $           � � C 7       �����&        x     ��  ��k       ���� � ������������+         ����
  % &           � � F :       �����'  �      x     ��  ��k       ���� � ������������+         ����
  ' (           � � I =       ����F(  �   	   x     ��  ��k       ���� � ������������+         ����
  ) *           � � L @       �����(  �      x     ��  ��k       ���� � ������������+         ����
  + ,           � � O C       �����)  �#      x	     ��  ��k       ���� � ������������+          ��              � � 4 ( P     �����!  ��        �       �     l        ���� � ������������,          ��              � � 7 + P     ����~"  r�        �      �     l        ���� � ������������,          ��              � � : . P     ����2#  ^�        �      �     l        ���� � ������������,          ��              � � = 1 P     �����#  J�        �      �     l        ���� � ������������,          ��    !           � � @ 4 P     �����$  6        �      �     l        ���� � ������������,          ��  # $           � � C 7 P     ����N%  "       �      �     l        ���� � ������������,          ��  % &           � � F : P     ����&  
       �      �     l        ���� � ������������,          ��  ' (           � � I = P     �����&  �       �      �     l        ���� � ������������,          ��  ) *           � � L @ P     ����j'  �       �      �     l        ���� � ������������,          ��  + ,           � � O C P     ����(  �       � 	     �     l        ���� � ������������,         ����              � � 4 (       ����
(  F      �      ��  ��m        ���� � ������������-         ����              � � 7 +       �����(  2      �     ��  ��m        ���� � ������������-         ����              � � : .       ����r)  "      �     ��  ��m        ���� � ������������-         ����               � � = 1       ����&*  
'      �     ��  ��m       ���� � ������������-         ����  ! "           � � @ 4       �����*  �+      �     ��  ��m       ���� � ������������-         ����  $ %           � � C 7       �����+  �0      �     ��  ��m       ���� � ������������-         ����  & '           � � F :       ����B,  �5      �     ��  ��m       ���� � ������������-         ����  ( )           � � I =       �����,  �:   	   �     ��  ��m       ���� � ������������-         ����  * +           � � L @       �����-  �?      �     ��  ��m       ���� � ������������-         ����  , -           � � O C       ����^.  �D      �	     ��  ��m       ���� � ������������-         ����	              � � 4 (       �����$  f            ��  ��n        ���� � ������������.         ����	              � � 7 +       �����%  R           ��  ��n        ���� � ������������.         ����	              � � : .       ����R&  >           ��  ��n        ���� � ������������.         ����	              � � = 1       ����'  *           ��  ��n       ���� � ������������.         ����	               � � @ 4       �����'             ��  ��n       ���� � ������������.         ����	  " #           � � C 7       ����n(             ��  ��n       ���� � ������������.         ����	  $ %           � � F :       ����")  �           ��  ��n       ���� � ������������.         ����	  & '           � � I =       �����)  �$   	        ��  ��n       ���� � ������������.         ����	  ( )           � � L @       �����*  �)           ��  ��n       ���� � ������������.         ����	  * +           � � O C       ����>+  �.      	     ��  ��n       ���� � ������������.         ����              � � 4 (       ����z&  V      ,      ��  ��o        ���� � ������������/         ����              � � 7 +       ����.'  B      ,     ��  ��o        ���� � ������������/         ����              � � : .       �����'  .      ,     ��  ��o        ���� � ������������/         ����               � � = 1       �����(        ,     ��  ��o       ���� � ������������/         ����  ! "           � � @ 4       ����J)  !      ,     ��  ��o       ���� � ������������/         ����  $ %           � � C 7       �����)  �%      ,     ��  ��o       ���� � ������������/         ����  & '           � � F :       �����*  �*      ,     ��  ��o       ���� � ������������/         ����  ( )           � � I =       ����f+  �/   	   ,     ��  ��o       ���� � ������������/         ����  * +           � � L @       ����,  �4      ,     ��  ��o       ���� � ������������/         ����  , -           � � O C       �����,  �9      ,	     ��  ��o       ���� � ������������/         ����              � � : .       �  #  �      l        ��p        ���� � �����  �  0         ����              � � > 2       �  �#  �      l       ��p        ���� � �����  �  0         ����               � � B 6       �  �$  &      l       ��p        ���� � �����  �  0         ����   ! "          � � F :         �%  �,      l       ��p       ���� � �����  �  0         ����   # $          � � J >         f&  03      l       ��p       ���� � �����  �  0         ����   % &          � � N B       #  8'  �9   	   l       ��p       ���� � �����  �  0         ����   ( )          � � R F       4  
(  P@      l       ��p       ���� � �����  �  0         ����   * +          � � V J       D  �(  �F      l       ��p       ���� � �����  �  0         ����   , -          � � Z N       U  �)  pM      l       ��p       ���� � �����  �  0         ����   . /          � � ^ R       f  �*   T      l	       ��p       ���� � �����  �  0         ����             � � : .       �  �   0      :        ��q        ���� � �����  �  1         ����             � � > 2       �  �!  �      :       ��q        ���� � �����  �  1         ����              � � B 6       �  j"  P      :       ��q        ���� � �����  �  1         ����  ! "          � � F :       �  <#  �      :       ��q       ���� � �����  �  1         ����  # $          � � J >       �  $  p       :       ��q       ���� � �����  �  1         ����  % &          � � N B       �  �$   '   	   :       ��q       ���� � �����  �  1         ����  ( )          � � R F         �%  �-      :       ��q       ���� � �����  �  1         ����  * +          � � V J         �&   4      :       ��q       ���� � �����  �  1         ����  , -          � � Z N       %  V'  �:      :       ��q       ���� � �����  �  1         ����  . /          � � ^ R       6  ((  @A      :	       ��q       ���� � �����  �  1         ����             � � : .       �  *!  P	      �        ��r        ���� � �����  �  2         ����             � � > 2       �  �!  �      �       ��r        ���� � �����  �  2         ����              � � B 6       �  �"  p      �       ��r        ���� � �����  �  2         ����  ! "          � � F :       �  �#         �       ��r       ���� � �����  �  2         ����  # $          � � J >       �  r$  �#      �       ��r       ���� � �����  �  2         ����  % &          � � N B       �  D%   *   	   �       ��r       ���� � �����  �  2         ����  ( )          � � R F         &  �0      �       ��r       ���� � �����  �  2         ����  * +          � � V J         �&  @7      �       ��r       ���� � �����  �  2         ����  , -          � � Z N       -  �'  �=      �       ��r       ���� � �����  �  2         ����  . /          � � ^ R       >  �(  `D      �	       ��r       ���� � �����  �  2         ����             � � : .       /  �'  p>      �        ��s        ���� � �����  �  3         ����             � � > 2       @  �(   E      �       ��s        ���� � �����  �  3         ����              � � B 6       P  r)  �K      �       ��s        ���� � �����  �  3         ����  ! "          � � F :       a  D*   R      �       ��s       ���� � �����  �  3         ����  # $          � � J >       r  +  �X      �       ��s       ���� � �����  �  3         ����  % &          � � N B       �  �+  @_   	   �       ��s       ���� � �����  �  3         ����  ( )          � � R F       �  �,  �e      �       ��s       ���� � �����  �  3         ����  * +          � � V J       �  �-  `l      �       ��s       ���� � �����  �  3         ����  , -          � � Z N       �  ^.  �r      �       ��s       ���� � �����  �  3         ����  . /          � � ^ R       �  0/  �y      �	       ��s       ���� � �����  �  3         ����             � � : .       �  �$  p%      l        ��t        ���� � �����  �  4         ����             � � > 2          �%   ,      l       ��t        ���� � �����  �  4         ����    !          � � B 6         R&  �2      l       ��t        ���� � �����  �  4         ����  " #          � � F :       !  $'   9      l       ��t       ���� � �����  �  4         ����  $ %          � � J >       2  �'  �?      l       ��t       ���� � �����  �  4         ����  & '          � � N B       C  �(  @F   	   l       ��t       ���� � �����  �  4         ����  ) *          � � R F       T  �)  �L      l       ��t       ���� � �����  �  4         ����  + ,          � � V J       d  l*  `S      l       ��t       ���� � �����  �  4         ����  - .          � � Z N       u  >+  �Y      l       ��t       ���� � �����  �  4         ����  / 0          � � ^ R       �  ,  �`      l	       ��t       ���� � �����  �  4         ����             � � : .         >&  �1              ��u        ���� � �����  �  5         ����              � � > 2          '  �8             ��u        ���� � �����  �  5         ����  ! "          � � B 6       0  �'  ?             ��u        ���� � �����  �  5         ����  # $          � � F :       A  �(  �E             ��u       ���� � �����  �  5         ����  % &          � � J >       R  �)  0L             ��u       ���� � �����  �  5         ����  ' (          � � N B       c  X*  �R   	          ��u       ���� � �����  �  5         ����  * +          � � R F       t  *+  PY             ��u       ���� � �����  �  5         ����  , -          � � V J       �  �+  �_             ��u       ���� � �����  �  5         ����  . /          � � Z N       �  �,  pf             ��u       ���� � �����  �  5         ����  0 1          � � ^ R       �  �-   m      	       ��u       ���� � �����  �  5         ����              � � : .       �����!  �      �      ��  ��v        ���� � �����  �  6         ����               � � > 2       �����"         �     ��  ��v        ���� � �����  �  6         ����  ! "           � � B 6       �����#  �      �     ��  ��v        ���� � �����  �  6         ����  # $           � � F :       ����h$  @#      �     ��  ��v       ���� � �����  �  6         ����  % &           � � J >       ����:%  �)      �     ��  ��v       ���� � �����  �  6         ����  ' (           � � N B       ����&  `0   	   �     ��  ��v       ���� � �����  �  6         ����  * +           � � R F       �����&  �6      �     ��  ��v       ���� � �����  �  6         ����  , -           � � V J       �����'  �=      �     ��  ��v       ���� � �����  �  6         ����  . /           � � Z N       �����(  D      �     ��  ��v       ���� � �����  �  6         ����  0 1           � � ^ R       ����T)  �J      �	     ��  ��v       ���� � �����  �  6         ����
              � � : .       ����~,  �c      y      ��  ��w        ���� � �����  �  7         ����
              � � > 2       ����P-  �j      y     ��  ��w        ���� � �����  �  7         ����
    !           � � B 6       ����".  q      y     ��  ��w        ���� � �����  �  7         ����
  " #           � � F :       �����.  �w      y     ��  ��w       ���� � �����  �  7         ����
  $ %           � � J >       �����/  0~      y     ��  ��w       ���� � �����  �  7         ����
  & '           � � N B       �����0  ��   	   y     ��  ��w       ���� � �����  �  7         ����
  ) *           � � R F       ����j1  P�      y     ��  ��w       ���� � �����  �  7         ����
  + ,           � � V J       ����<2  ��      y     ��  ��w       ���� � �����  �  7         ����
  - .           � � Z N       ����3  p�      y     ��  ��w       ���� � �����  �  7         ����
  / 0           � � ^ R       �����3   �      y	     ��  ��w       ���� � �����  �  7          ��              � � : . Z     �����*  pW       �       �     x        ���� � �����  �  8          ��              � � > 2 Z     �����+   ^       �      �     x        ���� � �����  �  8          ��    !           � � B 6 Z     �����,  �d       �      �     x        ���� � �����  �  8          ��  " #           � � F : Z     ����d-   k       �      �     x        ���� � �����  �  8          ��  $ %           � � J > Z     ����6.  �q       �      �     x        ���� � �����  �  8          ��  & '           � � N B Z     ����/  @x       �      �     x        ���� � �����  �  8          ��  ) *           � � R F Z     �����/  �~       �      �     x        ���� � �����  �  8          ��  + ,           � � V J Z     �����0  `�       �      �     x        ���� � �����  �  8          ��  - .           � � Z N Z     ����~1  ��       �      �     x        ���� � �����  �  8          ��  / 0           � � ^ R Z     ����P2  ��       � 	     �     x        ���� � �����  �  8         ����              � � : .       ����.1  p�      �      ��  ��y        ���� � �����  �  9         ����               � � > 2       ���� 2   �      �     ��  ��y        ���� � �����  �  9         ����  ! "           � � B 6       �����2  ��      �     ��  ��y        ���� � �����  �  9         ����  # $           � � F :       �����3   �      �     ��  ��y       ���� � �����  �  9         ����  % &           � � J >       ����v4  ��      �     ��  ��y       ���� � �����  �  9         ����  ' (           � � N B       ����H5  @�   	   �     ��  ��y       ���� � �����  �  9         ����  * +           � � R F       ����6  а      �     ��  ��y       ���� � �����  �  9         ����  , -           � � V J       �����6  `�      �     ��  ��y       ���� � �����  �  9         ����  . /           � � Z N       �����7  �      �     ��  ��y       ���� � �����  �  9         ����  0 1           � � ^ R       �����8  ��      �	     ��  ��y       ���� � �����  �  9         ����	              � � : .       ����.  pp            ��  ��z        ���� � �����  �  :         ����	              � � > 2       �����.   w           ��  ��z        ���� � �����  �  :         ����	               � � B 6       �����/  �}           ��  ��z        ���� � �����  �  :         ����	  ! "           � � F :       �����0   �           ��  ��z       ���� � �����  �  :         ����	  # $           � � J >       ����V1  ��           ��  ��z       ���� � �����  �  :         ����	  % &           � � N B       ����(2  @�   	        ��  ��z       ���� � �����  �  :         ����	  ( )           � � R F       �����2  З           ��  ��z       ���� � �����  �  :         ����	  * +           � � V J       �����3  `�           ��  ��z       ���� � �����  �  :         ����	  , -           � � Z N       �����4  �           ��  ��z       ���� � �����  �  :         ����	  . /           � � ^ R       ����p5  ��      	     ��  ��z       ���� � �����  �  :         ����              � � : .       �����/  �|      -      ��  ��{        ���� � �����  �  ;         ����               � � > 2       ����p0  ��      -     ��  ��{        ���� � �����  �  ;         ����  ! "           � � B 6       ����B1  �      -     ��  ��{        ���� � �����  �  ;         ����  # $           � � F :       ����2  ��      -     ��  ��{       ���� � �����  �  ;         ����  % &           � � J >       �����2  0�      -     ��  ��{       ���� � �����  �  ;         ����  ' (           � � N B       �����3  ��   	   -     ��  ��{       ���� � �����  �  ;         ����  * +           � � R F       �����4  P�      -     ��  ��{       ���� � �����  �  ;         ����  , -           � � V J       ����\5  �      -     ��  ��{       ���� � �����  �  ;         ����  . /           � � Z N       ����.6  p�      -     ��  ��{       ���� � �����  �  ;         ����  0 1           � � ^ R       ���� 7   �      -	     ��  ��{       ���� � �����  �  ;         ����  ' (            d �         2   `	  �        �      �   |        ����c   ������������<         ����  ) *            g �         0   ~	  �        �     �   |        ����c   ������������<         ����  + ,            j �         1   �	  8        �     �   |        ����c   ������������<         ����  - .            m �         1   �	  t        �     �   |       ����c   ������������<         ����  / 0            p �         2   �	  �        �     �   |       ����c   ������������<         ����  1 2            s �         3   �	  �        �     �   |       ����c   ������������<         ����  3 4            v �         3   
  (        �     �   |       ����c   ������������<         ����  5 6            y �         4   2
  d        �     �   |       ����c   ������������<         ����  7 8            | �         4   P
  �        �     �   |       ����c   ������������<         ����  9 :             �         5   n
  �        �	     �   |       ����c   ������������<         ����               � � J >         �-  �      m        ��}        ���� � �����  �  =         ����   ! "          � � N B       4  �.  x�      m       ��}        ���� � �����  �  =         ����   # $          � � R F       J  �/  �      m       ��}        ���� � �����  �  =         ����   % &          � � V J       _  �0  X�   	   m       ��}       ���� � �����  �  =         ����   ' (          � � Z N       u  �1  Ƚ      m       ��}       ���� � �����  �  =         ����   ) *          � � ^ R       �  x2  8�      m       ��}       ���� � �����  �  =         ����   , -          � � b V       �  h3  ��      m       ��}       ���� � �����  �  =         ����   . /          � � f Z       �  X4  �      m       ��}       ���� � �����  �  =         ����   0 1          � � j ^       �  H5  ��      m       ��}       ���� � �����  �  =         ����   2 3          � � n b       �  86  ��      m	       ��}       ���� � -  �  �  =         ����              � � J >       �  p+  ��      ;        ��~        ���� � �����  �  >         ����  ! "          � � N B       �  `,  `�      ;       ��~        ���� � �����  �  >         ����  # $          � � R F         P-  З      ;       ��~        ���� � �����  �  >         ����  % &          � � V J       )  @.  @�   	   ;       ��~       ���� � �����  �  >         ����  ' (          � � Z N       ?  0/  ��      ;       ��~       ���� � �����  �  >         ����  ) *          � � ^ R       T   0   �      ;       ��~       ���� � �����  �  >         ����  , -          � � b V       j  1  ��      ;       ��~       ���� � �����  �  >         ����  . /          � � f Z       �   2   �      ;       ��~       ���� � �����  �  >         ����  0 1          � � j ^       �  �2  p�      ;       ��~       ���� � �����  �  >         ����  2 3          � � n b       �  �3  ��      ;	       ��~       ���� � -  �  �  >         ����              � � J >       �  �+  t�      �        ��        ���� � �����  �  ?         ����  ! "          � � N B         �,  �      �       ��        ���� � �����  �  ?         ����  # $          � � R F         �-  T�      �       ��        ���� � �����  �  ?         ����  % &          � � V J       2  �.  ģ   	   �       ��       ���� � �����  �  ?         ����  ' (          � � Z N       H  �/  4�      �       ��       ���� � �����  �  ?         ����  ) *          � � ^ R       ]  �0  ��      �       ��       ���� � �����  �  ?         ����  , -          � � b V       s  t1  �      �       ��       ���� � �����  �  ?         ����  . /          � � f Z       �  d2  ��      �       ��       ���� � �����  �  ?         ����  0 1          � � j ^       �  T3  ��      �       ��       ���� � �����  �  ?         ����  2 3          � � n b       �  D4  d�      �	       ��       ���� � -  �  �  ?         ����              � � J >       �  x2  8�      �        ���        ���� � �����  �  @         ����  ! "          � � N B       �  h3  ��      �       ���        ���� � �����  �  @         ����  # $          � � R F       �  X4  �      �       ���        ���� � �����  �  @         ����  % &          � � V J       �  H5  ��   	   �       ���       ���� � �����  �  @         ����  ' (          � � Z N       �  86  ��      �       ���       ���� � �����  �  @         ����  ) *          � � ^ R       �  (7  h�      �       ���       ���� � �����  �  @         ����  , -          � � b V         8  ��      �       ���       ���� � �����  �  @         ����  . /          � � f Z       "  9  H      �       ���       ���� � �����  �  @         ����  0 1          � � j ^       7  �9  �	      �       ���       ���� � �����  �  @         ����  2 3          � � n b       M  �:  (      �	       ���       ���� � -  �  �  @         ����    !          � � J >       B  X/  �      m        ���        ���� � �����  �  A         ����  " #          � � N B       X  H0  ��      m       ���        ���� � �����  �  A         ����  $ %          � � R F       n  81  ��      m       ���        ���� � �����  �  A         ����  & '          � � V J       �  (2  h�   	   m       ���       ���� � �����  �  A         ����  ( )          � � Z N       �  3  ��      m       ���       ���� � �����  �  A         ����  * +          � � ^ R       �  4  H�      m       ���       ���� � �����  �  A         ����  - .          � � b V       �  �4  ��      m       ���       ���� � �����  �  A         ����  / 0          � � f Z       �  �5  (�      m       ���       ���� � �����  �  A         ����  1 2          � � j ^       �  �6  ��      m       ���       ���� � �����  �  A         ����  3 4          � � n b         �7  �      m	       ���       ���� � -  �  �  A         ����  ! "          � � J >       f  �0  (�              ���        ���� � �����  �  B         ����  # $          � � N B       |  �1  ��             ���        ���� � �����  �  B         ����  % &          � � R F       �  �2  �             ���        ���� � �����  �  B         ����  ' (          � � V J       �  �3  x�   	          ���       ���� � �����  �  B         ����  ) *          � � Z N       �  �4  ��             ���       ���� � �����  �  B         ����  + ,          � � ^ R       �  �5  X�             ���       ���� � �����  �  B         ����  . /          � � b V       �  �6  ��             ���       ���� � �����  �  B         ����  0 1          � � f Z       �  x7  8�             ���       ���� � �����  �  B         ����  2 3          � j ^         h8  ��             ���       ���� � �����  �  B         ����  4 5          � 	n b       )  X9        	       ���       ���� � -  �  �  B         ����  ! "           � � J >       �����,  |�      �      ��  ���        ���� � �����  �  C         ����  # $           � � N B       �����-  �      �     ��  ���        ���� � �����  �  C         ����  % &           � � R F       ����|.  \�      �     ��  ���        ���� � �����  �  C         ����  ' (           � � V J       ����l/  ̪   	   �     ��  ���       ���� � �����  �  C         ����  ) *           � � Z N       ����\0  <�      �     ��  ���       ���� � �����  �  C         ����  + ,           � � ^ R       ����L1  ��      �     ��  ���       ���� � �����  �  C         ����  . /           � � b V       ����<2  �      �     ��  ���       ���� � �����  �  C         ����  0 1           � � f Z       ����,3  ��      �     ��  ���       ���� � �����  �  C         ����  2 3           �  j ^       ����4  ��      �     ��  ���       ���� � �����  �  C         ����  4 5           � n b       ����5  l�      �	     ��  ���       ���� � �����  �  C         ����
    !           � � J >       ����(7  h�      z      ��  ���        ���� � �����  �  D         ����
  " #           � � N B       ����8  ��      z     ��  ���        ���� � �����  �  D         ����
  $ %           � � R F       ����9  H      z     ��  ���        ���� � �����  �  D         ����
  & '           � � V J       �����9  �	   	   z     ��  ���       ���� � �����  �  D         ����
  ( )           � � Z N       �����:  (      z     ��  ���       ���� � �����  �  D         ����
  * +           � � ^ R       �����;  �      z     ��  ���       ���� � �����  �  D         ����
  - .           � � b V       �����<  #      z     ��  ���       ���� � �����  �  D         ����
  / 0           � � f Z       �����=  x+      z     ��  ���       ���� � �����  �  D         ����
  1 2           � � j ^       �����>  �3      z     ��  ���       ���� � �����  �  D         ����
  3 4           � � n b       �����?  X<      z	     ��  ���       ���� � �����  �  D          ��    !           � � J > d     �����5  X�       �       �     �        ���� � �����  �  E          ��  " #           � � N B d     �����6  ��       �      �     �        ���� � �����  �  E          ��  $ %           � � R F d     ����x7  8�       �      �     �        ���� � �����  �  E          ��  & '           � � V J d     ����h8  ��       �      �     �        ���� � �����  �  E          ��  ( )           � � Z N d     ����X9         �      �     �        ���� � �����  �  E          ��  * +           � � ^ R d     ����H:  �       �      �     �        ���� � �����  �  E          ��  - .           � � b V d     ����8;  �       �      �     �        ���� � �����  �  E          ��  / 0           � � f Z d     ����(<  h       �      �     �        ���� � �����  �  E          ��  1 2           � j ^ d     ����=  �%       �      �     �        ���� � �����  �  E          ��  3 4           � 
n b d     ����>  H.       � 	     �     �        ���� � �����  �  E         ����  ! "           � � J >       �����;  �      �      ��  ���        ���� � �����  �  F         ����  # $           � � N B       �����<  #      �     ��  ���        ���� � �����  �  F         ����  % &           � � R F       �����=  x+      �     ��  ���        ���� � �����  �  F         ����  ' (           � � V J       �����>  �3   	   �     ��  ���       ���� � �����  �  F         ����  ) *           � � Z N       �����?  X<      �     ��  ���       ���� � �����  �  F         ����  + ,           � � ^ R       �����@  �D      �     ��  ���       ���� � �����  �  F         ����  . /           � � b V       ����xA  8M      �     ��  ���       ���� � �����  �  F         ����  0 1           � f Z       ����hB  �U      �     ��  ���       ���� � �����  �  F         ����  2 3           � 
j ^       ����XC  ^      �     ��  ���       ���� � �����  �  F         ����  4 5           � n b       ����HD  �f      �	     ��  ���       ���� � �����  �  F         ����	               � � J >       �����8  x�             ��  ���        ���� � �����  �  G         ����	  ! "           � � N B       �����9  �            ��  ���        ���� � �����  �  G         ����	  # $           � � R F       �����:  X            ��  ���        ���� � �����  �  G         ����	  % &           � � V J       �����;  �   	         ��  ���       ���� � �����  �  G         ����	  ' (           � � Z N       ����x<  8             ��  ���       ���� � �����  �  G         ����	  ) *           � � ^ R       ����h=  �(            ��  ���       ���� � �����  �  G         ����	  , -           � � b V       ����X>  1            ��  ���       ���� � �����  �  G         ����	  . /           � � f Z       ����H?  �9            ��  ���       ���� � �����  �  G         ����	  0 1           � � j ^       ����8@  �A            ��  ���       ���� � �����  �  G         ����	  2 3           � � n b       ����(A  hJ       	     ��  ���       ���� � �����  �  G         ����  ! "           � � J >       ����H:  �      .      ��  ���        ���� � �����  �  H         ����  # $           � � N B       ����8;  �      .     ��  ���        ���� � �����  �  H         ����  % &           � � R F       ����(<  h      .     ��  ���        ���� � �����  �  H         ����  ' (           � � V J       ����=  �%   	   .     ��  ���       ���� � �����  �  H         ����  ) *           � � Z N       ����>  H.      .     ��  ���       ���� � �����  �  H         ����  + ,           � � ^ R       �����>  �6      .     ��  ���       ���� � �����  �  H         ����  . /           � � b V       �����?  (?      .     ��  ���       ���� � �����  �  H         ����  0 1           � f Z       �����@  �G      .     ��  ���       ���� � �����  �  H         ����  2 3           � j ^       �����A  P      .     ��  ���       ���� � �����  �  H         ����  4 5           � n b       �����B  xX      .	     ��  ���       ���� � �����  �  H         ����   # $          � � Y M       �  �9  �C      n      	  ���        ����	 � �����  �  I         ����   % &          � � ] Q       �  ;  <N   
   n     	  ���        ����	 � �����  �  I         ����   ' (          � � a U         <  �X      n     	  ���        ����	 � �����  �  I         ����   ) *          � � e Y         "=  Tc      n     	  ���       ����	 � �����  �  I         ����   + ,          �  i ]       8  0>  �m      n     	  ���       ����	 � �����  �  I         ����   - .          � m a       S  >?  lx      n     	  ���       ����	 � �����  �  I         ����   0 1          � q e       n  L@  ��      n     	  ���       ����	 � �����  �  I         ����   2 3          u i       �  ZA  ��      n     	  ���       ����	 � �����  �  I         ����   4 5          
y m       �  hB  �       n     	  ���       ����	 � �����  �  I         ����   6 7          } q       �  vC  ��   ��  n	     	  ���       ����	 � 7  �  �  I         ����  # $          � � Y M       �  �7  @,      <      	  ���        ����	 � �����  �  J         ����  % &          � � ] Q       �  �8  �6   
   <     	  ���        ����	 � �����  �  J         ����  ' (          � � a U       �  �9  XA      <     	  ���        ����	 � �����  �  J         ����  ) *          � � e Y       �  �:  �K      <     	  ���       ����	 � �����  �  J         ����  + ,          � � i ]       �  �;  pV      <     	  ���       ����	 � �����  �  J         ����  - .          � m a         �<  �`      <     	  ���       ����	 � �����  �  J         ����  0 1          � q e       2  �=  �k      <     	  ���       ����	 � �����  �  J         ����  2 3          u i       M  ?  v      <     	  ���       ����	 � �����  �  J         ����  4 5          
y m       h  @  ��       <     	  ���       ����	 � �����  �  J         ����  6 7          } q       �  A  ,�   ��  <	     	  ���       ����	 � 7  �  �  J         ����  # $          � � Y M       �  8  (0      �      	  ���        ����	 � �����  �  K         ����  % &          � � ] Q       �  9  �:   
   �     	  ���        ����	 � �����  �  K         ����  ' (          � � a U       �   :  @E      �     	  ���        ����	 � �����  �  K         ����  ) *          � � e Y       �  .;  �O      �     	  ���       ����	 � �����  �  K         ����  + ,          � � i ]         <<  XZ      �     	  ���       ����	 � �����  �  K         ����  - .          � � m a       !  J=  �d      �     	  ���       ����	 � �����  �  K         ����  0 1          � q e       <  X>  po      �     	  ���       ����	 � �����  �  K         ����  2 3          u i       W  f?  �y      �     	  ���       ����	 � �����  �  K         ����  4 5          
y m       r  t@  ��       �     	  ���       ����	 � �����  �  K         ����  6 7          } q       �  �A  �   ��  �	     	  ���       ����	 � 7  �  �  K         ����  # $          � � Y M       D  �>  �r      �      	  ���        ����	 � �����  �  L         ����  % &          � � ] Q       _  �?  }   
   �     	  ���        ����	 � �����  �  L         ����  ' (          � � a U       z  �@  ��      �     	  ���        ����	 � �����  �  L         ����  ) *          � � e Y       �  �A  4�      �     	  ���       ����	 � �����  �  L         ����  + ,          � � i ]       �  �B  ��      �     	  ���       ����	 � �����  �  L         ����  - .          � � m a       �  �C  L�      �     	  ���       ����	 � �����  �  L         ����  0 1          � � q e       �  �D  ر      �     	  ���       ����	 � �����  �  L         ����  2 3          u i         
F  d�      �     	  ���       ����	 � �����  �  L         ����  4 5          
y m         G  ��       �     	  ���       ����	 � �����  �  L         ����  6 7          } q       7  &H  |�   ��  �	     	  ���       ����	 � 7  �  �  L         ����  $ %          � � Y M       �  �;  PS      n      	  ���        ����	 � �����  �  M         ����  & '          � � ] Q         �<  �]   
   n     	  ���        ����	 � �����  �  M         ����  ( )          � � a U       *  �=  hh      n     	  ���        ����	 � �����  �  M         ����  * +          � � e Y       E  �>  �r      n     	  ���       ����	 � �����  �  M         ����  , -          � � i ]       `  �?  �}      n     	  ���       ����	 � �����  �  M         ����  . /          � � m a       {  �@  �      n     	  ���       ����	 � �����  �  M         ����  1 2          � q e       �  �A  ��      n     	  ���       ����	 � �����  �  M         ����  3 4          	u i       �  �B  $�      n     	  ���       ����	 � �����  �  M         ����  5 6          
y m       �  �C  ��       n     	  ���       ����	 � �����  �  M         ����  7 8          } q       �  E  <�   ��  n	     	  ���       ����	 � 7  �  �  M         ����  % &          � � Y M         =  �b              ���        ����	 � �����  �  N         ����  ' (          � � ] Q       7  &>  |m   
          ���        ����	 � �����  �  N         ����  ) *          � � a U       R  4?  x             ���        ����	 � �����  �  N         ����  + ,          � e Y       m  B@  ��             ���       ����	 � �����  �  N         ����  - .          � 
i ]       �  PA   �             ���       ����	 � �����  �  N         ����  / 0          � m a       �  ^B  ��             ���       ����	 � �����  �  N         ����  2 3          � q e       �  lC  8�             ���       ����	 � �����  �  N         ����  4 5          u i       �  zD  Ĭ             ���       ����	 � �����  �  N         ����  6 7          
"y m       �  �E  P�              ���       ����	 � �����  �  N         ����  8 9          (} q         �F  ��   ��  	       ���       ����	 � 7  �  �  N         ����  % &           � � Y M       �����8  �7      �      ��  ���        ����	 � �����  �  O         ����  ' (           � � ] Q       �����9  �B   
   �     ��  ���        ����	 � �����  �  O         ����  ) *           � � a U       �����:  M      �     ��  ���        ����	 � �����  �  O         ����  + ,           � e Y       �����;  �W      �     ��  ���       ����	 � �����  �  O         ����  - .           � i ]       ����=  (b      �     ��  ���       ����	 � �����  �  O         ����  / 0           � m a       ����>  �l      �     ��  ���       ����	 � �����  �  O         ����  2 3           � q e       ���� ?  @w      �     ��  ���       ����	 � �����  �  O         ����  4 5           u i       ����.@  ́      �     ��  ���       ����	 � �����  �  O         ����  6 7           
y m       ����<A  X�       �     ��  ���       ����	 � �����  �  O         ����  8 9           %} q       ����JB  �   ��  �	     ��  ���       ����	 � �����  �  O         ����
  $ %           � � Y M       ����XC  p�      {      ��  ���        ����	 � �����  �  P         ����
  & '           � � ] Q       ����fD  ��   
   {     ��  ���        ����	 � �����  �  P         ����
  ( )           � � a U       ����tE  ��      {     ��  ���        ����	 � �����  �  P         ����
  * +           � � e Y       �����F  �      {     ��  ���       ����	 � �����  �  P         ����
  , -           � � i ]       �����G  ��      {     ��  ���       ����	 � �����  �  P         ����
  . /           � m a       �����H  ,�      {     ��  ���       ����	 � �����  �  P         ����
  1 2           � q e       �����I  ��      {     ��  ���       ����	 � �����  �  P         ����
  3 4           u i       �����J  D�      {     ��  ���       ����	 � �����  �  P         ����
  5 6           
y m       �����K  ��       {     ��  ���       ����	 � �����  �  P         ����
  7 8           } q       �����L  \    ��  {	     ��  ���       ����	 � �����  �  P          ��  $ %           � � Y M n     �����A  Б              �     �        ����	 � �����  �  Q          ��  & '           � � ] Q n     �����B  \�             �     �        ����	 � �����  �  Q          ��  ( )           � � a U n     �����C  �             �     �        ����	 � �����  �  Q          ��  * +           � e Y n     �����D  t�             �     �        ����	 � �����  �  Q          ��  , -           � i ] n     ���� F   �             �     �        ����	 � �����  �  Q          ��  . /           � m a n     ����G  ��             �     �        ����	 � �����  �  Q          ��  1 2           � q e n     ����H  �             �     �        ����	 � �����  �  Q          ��  3 4           u i n     ����*I  ��             �     �        ����	 � �����  �  Q          ��  5 6           
#y m n     ����8J  0�             �     �        ����	 � �����  �  Q          ��  7 8           )} q n     ����FK  ��        	     �     �        ����	 � �����  �  Q         ����  % &           � � Y M       ����H  P�      �      ��  ���        ����	 � �����  �  R         ����  ' (           � � ] Q       ����I  ��   
   �     ��  ���        ����	 � �����  �  R         ����  ) *           � a U       ����$J  h�      �     ��  ���        ����	 � �����  �  R         ����  + ,           � e Y       ����2K  ��      �     ��  ���       ����	 � �����  �  R         ����  - .           � i ]       ����@L  ��      �     ��  ���       ����	 � �����  �  R         ����  / 0           � m a       ����NM        �     ��  ���       ����	 � �����  �  R         ����  2 3           � q e       ����\N  �      �     ��  ���       ����	 � �����  �  R         ����  4 5           #u i       ����jO  $      �     ��  ���       ����	 � �����  �  R         ����  6 7           
)y m       ����xP  �$       �     ��  ���       ����	 � �����  �  R         ����  8 9           /} q       �����Q  </   ��  �	     ��  ���       ����	 � �����  �  R         ����	  # $           � � Y M       �����D  �      !      ��  ���        ����	 � �����  �  S         ����	  % &           � � ] Q       �����E  ��   
   !     ��  ���        ����	 � �����  �  S         ����	  ' (           � � a U       ����G  (�      !     ��  ���        ����	 � �����  �  S         ����	  ) *           � � e Y       ����H  ��      !     ��  ���       ����	 � �����  �  S         ����	  + ,           � � i ]       ���� I  @�      !     ��  ���       ����	 � �����  �  S         ����	  - .           � � m a       ����.J  ��      !     ��  ���       ����	 � �����  �  S         ����	  0 1           � q e       ����<K  X�      !     ��  ���       ����	 � �����  �  S         ����	  2 3           	u i       ����JL  ��      !     ��  ���       ����	 � �����  �  S         ����	  4 5           
y m       ����XM  p       !     ��  ���       ����	 � �����  �  S         ����	  6 7           } q       ����fN  �   ��  !	     ��  ���       ����	 � �����  �  S         ����  % &           � � Y M       ����xF  ��      /      ��  ���        ����	 � �����  �  T         ����  ' (           � � ] Q       �����G  <�   
   /     ��  ���        ����	 � �����  �  T         ����  ) *           � a U       �����H  ��      /     ��  ���        ����	 � �����  �  T         ����  + ,           � 	e Y       �����I  T�      /     ��  ���       ����	 � �����  �  T         ����  - .           � i ]       �����J  ��      /     ��  ���       ����	 � �����  �  T         ����  / 0           � m a       �����K  l�      /     ��  ���       ����	 � �����  �  T         ����  2 3           � q e       �����L  ��      /     ��  ���       ����	 � �����  �  T         ����  4 5           !u i       �����M  �
      /     ��  ���       ����	 � �����  �  T         ����  6 7           
'y m       �����N         /     ��  ���       ����	 � �����  �  T         ����  8 9           -} q       �����O  �   ��  /	     ��  ���       ����	 � �����  �  T         ����   ' (          � h \       �  �G  z   	   o      
  ���        ����
 � �����  �  U         ����   ) *           l `         �H  ^!      o     
  ���        ����
 � �����  �  U         ����   + ,          p d       $  J  B.      o     
  ���        ����
 � �����  �  U         ����   - .          t h       E  2K  &;      o     
  ���       ����
 � �����  �  U         ����   / 0          x l       f  ^L  
H      o     
  ���       ����
 � �����  �  U         ����   1 2          $| p       �  �M  �T      o     
  ���       ����
 � �����  �  U         ����   4 5          *� t       �  �N  �a      o     
  ���       ����
 � �����  �  U         ����   6 7          $0� x       �  �O  �n   ��  o     
  ���       ����
 � �����  �  U         ����   8 9          *6� |       �  Q  �{   ��  o     
  ���       ����
 � �����  �  U         ����   : ;          0<� �       	  :R  ~�   ��  o	     
  ���       ����
 7  �  �  U         ����  ' (          � h \       �  VE  ��   	   =      
  ���        ����
 � �����  �  V         ����  ) *           l `       �  �F  �      =     
  ���        ����
 � �����  �  V         ����  + ,          p d       �  �G  z      =     
  ���        ����
 � �����  �  V         ����  - .          t h         �H  ^!      =     
  ���       ����
 � �����  �  V         ����  / 0          x l       $  J  B.      =     
  ���       ����
 � �����  �  V         ����  1 2          #| p       E  2K  &;      =     
  ���       ����
 � �����  �  V         ����  4 5          )� t       f  ^L  
H      =     
  ���       ����
 � �����  �  V         ����  6 7          $/� x       �  �M  �T   ��  =     
  ���       ����
 � �����  �  V         ����  8 9          *5� |       �  �N  �a   ��  =     
  ���       ����
 � �����  �  V         ����  : ;          0;� �       �  �O  �n   ��  =	     
  ���       ����
 7  �  �  V         ����  ' (          � � h \       �  �E  ��   	   �      
  ���        ����
 � �����  �  W         ����  ) *           l `       �  �F  �      �     
  ���        ����
 � �����  �  W         ����  + ,          p d       �  H  �      �     
  ���        ����
 � �����  �  W         ����  - .          t h         >I  �%      �     
  ���       ����
 � �����  �  W         ����  / 0          x l       /  jJ  �2      �     
  ���       ����
 � �����  �  W         ����  1 2          | p       P  �K  r?      �     
  ���       ����
 � �����  �  W         ����  4 5           � t       q  �L  VL      �     
  ���       ����
 � �����  �  W         ����  6 7          $&� x       �  �M  :Y   ��  �     
  ���       ����
 � �����  �  W         ����  8 9          *,� |       �  O  f   ��  �     
  ���       ����
 � �����  �  W         ����  : ;          02� �       �  FP  s   ��  �	     
  ���       ����
 7  �  �  W         ����  ' (          � � h \       f  ^L  
H   	   �      
  ���        ����
 � �����  �  X         ����  ) *           � l `       �  �M  �T      �     
  ���        ����
 � �����  �  X         ����  + ,          p d       �  �N  �a      �     
  ���        ����
 � �����  �  X         ����  - .          t h       �  �O  �n      �     
  ���       ����
 � �����  �  X         ����  / 0          x l       �  Q  �{      �     
  ���       ����
 � �����  �  X         ����  1 2          | p       	  :R  ~�      �     
  ���       ����
 � �����  �  X         ����  4 5          � t       ,	  fS  b�      �     
  ���       ����
 � �����  �  X         ����  6 7          $#� x       M	  �T  F�   ��  �     
  ���       ����
 � �����  �  X         ����  8 9          *)� |       n	  �U  *�   ��  �     
  ���       ����
 � �����  �  X         ����  : ;          0/� �       �	  �V  �   ��  �	     
  ���       ����
 7  �  �  X         ����  ( )          � � h \         >I  �%   	   o      
  ���        ����
 � �����  �  Y         ����  * +           l `       /  jJ  �2      o     
  ���        ����
 � �����  �  Y         ����  , -          	p d       P  �K  r?      o     
  ���        ����
 � �����  �  Y         ����  . /          t h       q  �L  VL      o     
  ���       ����
 � �����  �  Y         ����  0 1          x l       �  �M  :Y      o     
  ���       ����
 � �����  �  Y         ����  2 3          | p       �  O  f      o     
  ���       ����
 � �����  �  Y         ����  5 6          !� t       �  FP  s      o     
  ���       ����
 � �����  �  Y         ����  7 8          $'� x       �  rQ  �   ��  o     
  ���       ����
 � �����  �  Y         ����  9 :          *-� |       	  �R  ʌ   ��  o     
  ���       ����
 � �����  �  Y         ����  ; <          03� �       7	  �S  ��   ��  o	     
  ���       ����
 7  �  �  Y         ����  ) *          � h \       :  �J  �6   	   	      	  ���        ����
 � �����  �  Z         ����  + ,           l `       [  �K  �C      	     	  ���        ����
 � �����  �  Z         ����  - .          p d       |  &M  �P      	     	  ���        ����
 � �����  �  Z         ����  / 0          "t h       �  RN  �]      	     	  ���       ����
 � �����  �  Z         ����  1 2          (x l       �  ~O  jj      	     	  ���       ����
 � �����  �  Z         ����  3 4          .| p       �  �P  Nw      	     	  ���       ����
 � �����  �  Z         ����  6 7          4� t        	  �Q  2�      	     	  ���       ����
 � �����  �  Z         ����  8 9          $:� x       !	  S  �   ��  	     	  ���       ����
 � �����  �  Z         ����  : ;          *@� |       B	  .T  ��   ��  	     	  ���       ����
 � �����  �  Z         ����  < =          0F� �       c	  ZU  ު   ��  		     	  ���       ����
 7  �  �  Z         ����  ) *           � h \       �����F  �   	   �      ��  ���        ����
 � �����  �  [         ����  + ,            l `       �����G  z      �     ��  ���        ����
 � �����  �  [         ����  - .           p d       �����H  ^!      �     ��  ���        ����
 � �����  �  [         ����  / 0           t h       ����J  B.      �     ��  ���       ����
 � �����  �  [         ����  1 2           %x l       ����2K  &;      �     ��  ���       ����
 � �����  �  [         ����  3 4           +| p       ����^L  
H      �     ��  ���       ����
 � �����  �  [         ����  6 7           1� t       �����M  �T      �     ��  ���       ����
 � �����  �  [         ����  8 9           $7� x       �����N  �a   ��  �     ��  ���       ����
 � �����  �  [         ����  : ;           *=� |       �����O  �n   ��  �     ��  ���       ����
 � �����  �  [         ����  < =           0C� �       ����Q  �{   ��  �	     ��  ���       ����
 �����  �  [         ����
  ( )           � h \       ����Q  �{   	   |      ��  ���        ����
 � �����  �  \         ����
  * +            l `       ����:R  ~�      |     ��  ���        ����
 � �����  �  \         ����
  , -           p d       ����fS  b�      |     ��  ���        ����
 � �����  �  \         ����
  . /           t h       �����T  F�      |     ��  ���       ����
 � �����  �  \         ����
  0 1           x l       �����U  *�      |     ��  ���       ����
 � �����  �  \         ����
  2 3           #| p       �����V  �      |     ��  ���       ����
 � �����  �  \         ����
  5 6           )� t       ����X  ��      |     ��  ���       ����
 � �����  �  \         ����
  7 8           $/� x       ����BY  ��   ��  |     ��  ���       ����
 � �����  �  \         ����
  9 :           *5� |       ����nZ  ��   ��  |     ��  ���       ����
 � �����  �  \         ����
  ; <           0;� �       �����[  ��   ��  |	     ��  ���       ����
 �����  �  \          ��  ( )           � h \ x     ����~O  jj             �     �        ����
 � �����  �  ]          ��  * +            l ` x     �����P  Nw            �     �        ����
 � �����  �  ]          ��  , -           p d x     �����Q  2�            �     �        ����
 � �����  �  ]          ��  . /           #t h x     ����S  �            �     �        ����
 � �����  �  ]          ��  0 1           )x l x     ����.T  ��            �     �        ����
 � �����  �  ]          ��  2 3           /| p x     ����ZU  ު            �     �        ����
 � �����  �  ]          ��  5 6           5� t x     �����V  ·            �     �        ����
 � �����  �  ]          ��  7 8           $;� x x     �����W  ��            �     �        ����
 � �����  �  ]          ��  9 :           *A� | x     �����X  ��            �     �        ����
 � �����  �  ]          ��  ; <           0G� � x     ����
Z  n�       	     �     �        ����
 �����  �  ]         ����  ) *           � h \       �����U  *�   	   �      ��  ���        ����
 � �����  �  ^         ����  + ,            l `       �����V  �      �     ��  ���        ����
 � �����  �  ^         ����  - .           #p d       ����X  ��      �     ��  ���        ����
 � �����  �  ^         ����  / 0           )t h       ����BY  ��      �     ��  ���       ����
 � �����  �  ^         ����  1 2           /x l       ����nZ  ��      �     ��  ���       ����
 � �����  �  ^         ����  3 4           5| p       �����[  ��      �     ��  ���       ����
 � �����  �  ^         ����  6 7           ;� t       �����\  ��      �     ��  ���       ����
 � �����  �  ^         ����  8 9           $A� x       �����]  f	   ��  �     ��  ���       ����
 � �����  �  ^         ����  : ;           *G� |       ����_  J   ��  �     ��  ���       ����
 � �����  �  ^         ����  < =           0M� �       ����J`  .#   ��  �	     ��  ���       ����
 �����  �  ^         ����	  ' (           � � h \       �����R  ʌ   	   "      ��  ���        ����
 � �����  �  _         ����	  ) *            l `       �����S  ��      "     ��  ���        ����
 � �����  �  _         ����	  + ,           	p d       �����T  ��      "     ��  ���        ����
 � �����  �  _         ����	  - .           t h       ����"V  v�      "     ��  ���       ����
 � �����  �  _         ����	  / 0           x l       ����NW  Z�      "     ��  ���       ����
 � �����  �  _         ����	  1 2           | p       ����zX  >�      "     ��  ���       ����
 � �����  �  _         ����	  4 5           !� t       �����Y  "�      "     ��  ���       ����
 � �����  �  _         ����	  6 7           $'� x       �����Z  �   ��  "     ��  ���       ����
 � �����  �  _         ����	  8 9           *-� |       �����[  ��   ��  "     ��  ���       ����
 � �����  �  _         ����	  : ;           03� �       ����*]  �    ��  "	     ��  ���       ����
 �����  �  _         ����  ) *           � h \       ����.T  ��   	   0      ��  ���        ����
 � �����  �  `         ����  + ,            l `       ����ZU  ު      0     ��  ���        ����
 � �����  �  `         ����  - .           !p d       �����V  ·      0     ��  ���        ����
 � �����  �  `         ����  / 0           't h       �����W  ��      0     ��  ���       ����
 � �����  �  `         ����  1 2           -x l       �����X  ��      0     ��  ���       ����
 � �����  �  `         ����  3 4           3| p       ����
Z  n�      0     ��  ���       ����
 � �����  �  `         ����  6 7           9� t       ����6[  R�      0     ��  ���       ����
 � �����  �  `         ����  8 9           $?� x       ����b\  6�   ��  0     ��  ���       ����
 � �����  �  `         ����  : ;           *E� |       �����]     ��  0     ��  ���       ����
 � �����  �  `         ����  < =           0K� �       �����^  �   ��  0	     ��  ���       ����
 �����  �  `         ����   + ,          #v j d     n
  �V  �      p        ���        ���� � �����  �  a         ����   - .           *{ o e     �
  4X  p"      p       ���        ���� � �����  �  a         ����   / 0          '1� t f     �
  ~Y  �1      p       ���        ���� � �����  �  a         ����   1 2          .8� y g     �
  �Z  `A      p       ���       ���� � �����  �  a         ����   3 4          5?� ~ h       \  �P      p       ���       ���� � �����  �  a         ����   5 6          <F� � i     4  \]  P`   ��  p       ���       ���� � �����  �  a         ����   8 9          CM� � j     [  �^  �o   ��  p       ���       ���� � �����  �  a         ����   : ;          JT� � k     �  �_  @   ��  p       ���       ���� � �����  �  a         ����   < =          Q[� � l     �  :a  ��   ��  p       ���       ���� �����  �  a         ����   > ?          Xb� � m     �  �b  0�   ��  p	       ���       ���� A  �  �  a         ����  + ,          "v j d     &
  �T  ��      >        ���        ���� � �����  �  b         ����  - .           ){ o e     M
  �U  P      >       ���        ���� � �����  �  b         ����  / 0          '0� t f     u
  &W  �      >       ���        ���� � �����  �  b         ����  1 2          .7� y g     �
  pX  @%      >       ���       ���� � �����  �  b         ����  3 4          5>� ~ h     �
  �Y  �4      >       ���       ���� � �����  �  b         ����  5 6          <E� � i     �
  [  0D   ��  >       ���       ���� � �����  �  b         ����  8 9          CL� � j       N\  �S   ��  >       ���       ���� � �����  �  b         ����  : ;          JS� � k     ;  �]   c   ��  >       ���       ���� � �����  �  b         ����  < =          QZ� � l     b  �^  �r   ��  >       ���       ���� �����  �  b         ����  > ?          Xa� � m     �  ,`  �   ��  >	       ���       ���� A  �  �  b         ����  + ,          v j d     2
  �T  ��      �        ���        ���� � �����  �  c         ����  - .            { o e     Y
  @V         �       ���        ���� � �����  �  c         ����  / 0          ''� t f     �
  �W  x      �       ���        ���� � �����  �  c         ����  1 2          ..� y g     �
  �X  �)      �       ���       ���� � �����  �  c         ����  3 4          55� ~ h     �
  Z  h9      �       ���       ���� � �����  �  c         ����  5 6          <<� � i     �
  h[  �H   ��  �       ���       ���� � �����  �  c         ����  8 9          CC� � j       �\  XX   ��  �       ���       ���� � �����  �  c         ����  : ;          JJ� � k     G  �]  �g   ��  �       ���       ���� � �����  �  c         ����  < =          QQ� � l     n  F_  Hw   ��  �       ���       ���� �����  �  c         ����  > ?          XX� � m     �  �`  ��   ��  �	       ���       ���� A  �  �  c         ����  + ,          v j d     �
  �[  8K      �        ���        ���� � �����  �  d         ����  - .           { o e     %  �\  �Z      �       ���        ���� � �����  �  d         ����  / 0          '$� t f     M  .^  (j      �       ���        ���� � �����  �  d         ����  1 2          .+� y g     t  x_  �y      �       ���       ���� � �����  �  d         ����  3 4          52� ~ h     �  �`  �      �       ���       ���� � �����  �  d         ����  5 6          <9� � i     �  b  ��   ��  �       ���       ���� � �����  �  d         ����  8 9          C@� � j     �  Vc  �   ��  �       ���       ���� � �����  �  d         ����  : ;          JG� � k       �d  ��   ��  �       ���       ���� � �����  �  d         ����  < =          QN� � l     :  �e  ��   ��  �       ���       ���� �����  �  d         ����  > ?          XU� � m     b  4g  p�   ��  �	       ���       ���� A  �  �  d         ����  , -          v j d     �
  zX  �%      p        ���        ���� � �����  �  e         ����  . /           !{ o e     �
  �Y  05      p       ���        ���� � �����  �  e         ����  0 1          '(� t f     �
  [  �D      p       ���        ���� � �����  �  e         ����  2 3          ./� y g       X\   T      p       ���       ���� � �����  �  e         ����  4 5          56� ~ h     <  �]  �c      p       ���       ���� � �����  �  e         ����  6 7          <=� � i     d  �^  s   ��  p       ���       ���� � �����  �  e         ����  9 :          CD� � j     �  6`  ��   ��  p       ���       ���� � �����  �  e         ����  ; <          JK� � k     �  �a   �   ��  p       ���       ���� � �����  �  e         ����  = >          QR� � l     �  �b  x�   ��  p       ���       ���� �����  �  e         ����  ? @          XY� � m       d  �   ��  p	       ���       ���� A  �  �  e         ����  - .          -v j d     �
  
Z  x8      
      
  ���        ���� � �����  �  f         ����  / 0           4{ o e     �
  T[  �G      
     
  ���        ���� � �����  �  f         ����  1 2          ';� t f       �\  hW      
     
  ���        ���� � �����  �  f         ����  3 4          .B� y g     D  �]  �f      
     
  ���       ���� � �����  �  f         ����  5 6          5I� ~ h     l  2_  Xv      
     
  ���       ���� � �����  �  f         ����  7 8          <P� � i     �  |`  Ѕ   ��  
     
  ���       ���� � �����  �  f         ����  : ;          CW� � j     �  �a  H�   ��  
     
  ���       ���� � �����  �  f         ����  < =          J^� � k     �  c  ��   ��  
     
  ���       ���� � �����  �  f         ����  > ?          Qe� � l     
  Zd  8�   ��  
     
  ���       ���� �����  �  f         ����  @ A          Xl� � m     2  �e  ��   ��  
	     
  ���       ���� A  �  �  f         ����  - .           *v j d     �����U  �      �      ��  ���        ���� � �����  �  g         ����  / 0            1{ o e     ����W  `      �     ��  ���        ���� � �����  �  g         ����  1 2           '8� t f     ����RX  �#      �     ��  ���        ���� � �����  �  g         ����  3 4           .?� y g     �����Y  P3      �     ��  ���       ���� � �����  �  g         ����  5 6           5F� ~ h     �����Z  �B      �     ��  ���       ���� � �����  �  g         ����  7 8           <M� � i     ����0\  @R   ��  �     ��  ���       ���� � �����  �  g         ����  : ;           CT� � j     ����z]  �a   ��  �     ��  ���       ���� � �����  �  g         ����  < =           J[� � k     �����^  0q   ��  �     ��  ���       ���� � �����  �  g         ����  > ?           Qb� � l     ����`  ��   ��  �     ��  ���       ���� �����  �  g         ����  @ A           Xi� � m     ����Xa   �   ��  �	     ��  ���       ���� �����  �  g         ����
  , -           "v j d     ����J`  x�      }      ��  ���        ���� � �����  �  h         ����
  . /            ){ o e     �����a  �      }     ��  ���        ���� � �����  �  h         ����
  0 1           '0� t f     �����b  h�      }     ��  ���        ���� � �����  �  h         ����
  2 3           .7� y g     ����(d  �      }     ��  ���       ���� � �����  �  h         ����
  4 5           5>� ~ h     ����re  X�      }     ��  ���       ���� � �����  �  h         ����
  6 7           <E� � i     �����f  ��   ��  }     ��  ���       ���� � �����  �  h         ����
  9 :           CL� � j     ����h  H�   ��  }     ��  ���       ���� � �����  �  h         ����
  ; <           JS� � k     ����Pi  ��   ��  }     ��  ���       ���� � �����  �  h         ����
  = >           QZ� � l     �����j  8�   ��  }     ��  ���       ���� �����  �  h         ����
  ? @           Xa� � m     �����k  �   ��  }	     ��  ���       ���� �����  �  h          ��  , -           .v j �     �����^  �p             �     �        ���� � �����  �  i          ��  . /            5{ o �     ����`  0�            �     �        ���� � �����  �  i          ��  0 1           '<� t �     ����Na  ��            �     �        ���� � �����  �  i          ��  2 3           .C� y �     �����b   �            �     �        ���� � �����  �  i          ��  4 5           5J� ~ �     �����c  ��            �     �        ���� � �����  �  i          ��  6 7           <Q� � �     ����,e  �            �     �        ���� � �����  �  i          ��  9 :           CX� � �     ����vf  ��            �     �        ���� � �����  �  i          ��  ; <           J_� � �     �����g   �            �     �        ���� � �����  �  i          ��  = >           Qf� � �     ����
i  x�            �     �        ���� �����  �  i          ��  ? @           Xm� � �     ����Tj  ��       	     �     �        ���� �����  �  i         ����  - .           4v j d     �����d  ��      �      ��  ���        ���� � �����  �  j         ����  / 0            ;{ o e     ����Df  0�      �     ��  ���        ���� � �����  �  j         ����  1 2           'B� t f     �����g  ��      �     ��  ���        ���� � �����  �  j         ����  3 4           .I� y g     �����h   �      �     ��  ���       ���� � �����  �  j         ����  5 6           5P� ~ h     ����"j  ��      �     ��  ���       ���� � �����  �  j         ����  7 8           <W� � i     ����lk  	   ��  �     ��  ���       ���� � �����  �  j         ����  : ;           C^� � j     �����l  �   ��  �     ��  ���       ���� � �����  �  j         ����  < =           Je� � k     ���� n   (   ��  �     ��  ���       ���� � �����  �  j         ����  > ?           Ql� � l     ����Jo  x7   ��  �     ��  ���       ���� �����  �  j         ����  @ A           Xs� � m     �����p  �F   ��  �	     ��  ���       ���� �����  �  j         ����	  + ,           v j d     �����a  8�      #      ��  ���        ���� � �����  �  k         ����	  - .            !{ o e     ����$c  ��      #     ��  ���        ���� � �����  �  k         ����	  / 0           '(� t f     ����nd  (�      #     ��  ���        ���� � �����  �  k         ����	  1 2           ./� y g     �����e  ��      #     ��  ���       ���� � �����  �  k         ����	  3 4           56� ~ h     ����g  �      #     ��  ���       ���� � �����  �  k         ����	  5 6           <=� � i     ����Lh  ��   ��  #     ��  ���       ���� � �����  �  k         ����	  8 9           CD� � j     �����i  �   ��  #     ��  ���       ���� � �����  �  k         ����	  : ;           JK� � k     �����j  �   ��  #     ��  ���       ���� � �����  �  k         ����	  < =           QR� � l     ����*l  �   ��  #     ��  ���       ���� �����  �  k         ����	  > ?           XY� � m     ����tm  p!   ��  #	     ��  ���       ���� �����  �  k         ����  - .           2v j d     ����jc  ��      1      ��  ���        ���� � �����  �  l         ����  / 0            9{ o e     �����d  p�      1     ��  ���        ���� � �����  �  l         ����  1 2           '@� t f     �����e  ��      1     ��  ���        ���� � �����  �  l         ����  3 4           .G� y g     ����Hg  `�      1     ��  ���       ���� � �����  �  l         ����  5 6           5N� ~ h     �����h  ��      1     ��  ���       ���� � �����  �  l         ����  7 8           <U� � i     �����i  P�   ��  1     ��  ���       ���� � �����  �  l         ����  : ;           C\� � j     ����&k  �   ��  1     ��  ���       ���� � �����  �  l         ����  < =           Jc� � k     ����pl  @   ��  1     ��  ���       ���� � �����  �  l         ����  > ?           Qj� � l     �����m  �$   ��  1     ��  ���       ���� �����  �  l         ����  @ A           Xq� � m     ����o  04   ��  1	     ��  ���       ���� �����  �  l         ����   / 0          AI� � n     z  �g  �C      q        ���        ���� � �����  �  m         ����   1 2          HP� � o     �  i  V      q       ���        ���� � �����  �  m         ����   3 4          OW� � p     �  |j  Lh      q       ���        ���� � �����  �  m         ����   5 6          V^� � q       �k  �z   ��  q       ���       ���� � �����  �  m         ����   7 8          ]e� � r     5  Lm  ܌   ��  q       ���       ���� � �����  �  m         ����   9 :          dl� � s     d  �n  $�   ��  q       ���       ���� � �����  �  m         ����   < =          ks� � t     �  p  l�   ��  q       ���       ����  �����  �  m         ����   > ?          rz� � u     �  �q  ��   ��  q       ���       ���� �����  �  m         ����   @ A          y�� � v     �  �r  ��   ��  q       ���       ���� �����  �  m         ����   B C          ��� � w       Tt  D�   ��  q	       ���       ���� A  �  �  m         ����  / 0          AH� � n     ,  Te  D%      ?        ���        ���� � �����  �  n         ����  1 2          HO� � o     [  �f  �7      ?       ���        ���� � �����  �  n         ����  3 4          OV� � p     �  $h  �I      ?       ���        ���� � �����  �  n         ����  5 6          V]� � q     �  �i  \   ��  ?       ���       ���� � �����  �  n         ����  7 8          ]d� � r     �  �j  dn   ��  ?       ���       ���� � �����  �  n         ����  9 :          dk� � s       \l  ��   ��  ?       ���       ���� � �����  �  n         ����  < =          kr� � t     E  �m  ��   ��  ?       ���       ����  �����  �  n         ����  > ?          ry� � u     s  ,o  <�   ��  ?       ���       ���� �����  �  n         ����  @ A          y�� � v     �  �p  ��   ��  ?       ���       ���� �����  �  n         ����  B C          ��� � w     �  �q  ��   ��  ?	       ���       ���� A  �  �  n         ����  / 0          A?� � n     9  �e  X*      �        ���        ���� � �����  �  o         ����  1 2          HF� � o     h   g  �<      �       ���        ���� � �����  �  o         ����  3 4          OM� � p     �  �h  �N      �       ���        ���� � �����  �  o         ����  5 6          VT� � q     �  �i  0a   ��  �       ���       ���� � �����  �  o         ����  7 8          ][� � r     �  Xk  xs   ��  �       ���       ���� � �����  �  o         ����  9 :          db� � s     #  �l  ��   ��  �       ���       ���� � �����  �  o         ����  < =          ki� � t     R  (n  �   ��  �       ���       ����  �����  �  o         ����  > ?          rp� � u     �  �o  P�   ��  �       ���       ���� �����  �  o         ����  @ A          yw� � v     �  �p  ��   ��  �       ���       ���� �����  �  o         ����  B C          �~� � w     �  `r  ��   ��  �	       ���       ���� A  �  �  o         ����  / 0          A<� � n       \l  ��      �        ���        ���� � �����  �  p         ����  1 2          HC� � o     E  �m  ��      �       ���        ���� � �����  �  p         ����  3 4          OJ� � p     s  ,o  <�      �       ���        ���� � �����  �  p         ����  5 6          VQ� � q     �  �p  ��   ��  �       ���       ���� � �����  �  p         ����  7 8          ]X� � r     �  �q  ��   ��  �       ���       ���� � �����  �  p         ����  9 :          d_� � s        ds  �   ��  �       ���       ���� � �����  �  p         ����  < =          kf� � t     /  �t  \�   ��  �       ���       ����  �����  �  p         ����  > ?          rm� � u     ]  4v  �    ��  �       ���       ���� �����  �  p         ����  @ A          yt� � v     �  �w  �   ��  �       ���       ���� �����  �  p         ����  B C          �{� � w     �  y  4%   ��  �	       ���       ���� A  �  �  p         ����  0 1          A@� � n     �  <i  X      q        ���        ���� � �����  �  q         ����  2 3          HG� � o     �  �j  Tj      q       ���        ���� � �����  �  q         ����  4 5          ON� � p       l  �|      q       ���        ���� � �����  �  q         ����  6 7          VU� � q     :  tm  �   ��  q       ���       ���� � �����  �  q         ����  8 9          ]\� � r     i  �n  ,�   ��  q       ���       ���� � �����  �  q         ����  : ;          dc� � s     �  Dp  t�   ��  q       ���       ���� � �����  �  q         ����  = >          kj� � t     �  �q  ��   ��  q       ���       ����  �����  �  q         ����  ? @          rq� � u     �  s  �   ��  q       ���       ���� �����  �  q         ����  A B          yx� � v     $  |t  L�   ��  q       ���       ���� �����  �  q         ����  C D          �� � w     S  �u  ��   ��  q	       ���       ���� A  �  �  q         ����  1 2          AS� � n     �  �j  \l              ���        ���� � �����  �  r         ����  3 4          HZ� � o       4l  �~             ���        ���� � �����  �  r         ����  5 6          Oa� � p     ?  �m  �             ���        ���� � �����  �  r         ����  7 8          Vh� � q     n  o  4�   ��         ���       ���� � �����  �  r         ����  9 :          ]o� � r     �  lp  |�   ��         ���       ���� � �����  �  r         ����  ; <          dv� � s     �  �q  ��   ��         ���       ���� � �����  �  r         ����  > ?          k}� � t     �  <s  �   ��         ���       ����  �����  �  r         ����  @ A          r�� � u     )  �t  T�   ��         ���       ���� �����  �  r         ����  B C          y�� � v     X  v  ��   ��         ���       ���� �����  �  r         ����  D E          ��� � w     �  tw  �   ��  	       ���       ���� A  �  �  r         ����  1 2           AP� � n     �����f  �4      �      ��  ���        ���� � �����  �  s         ����  3 4           HW� � o     �����g  �F      �     ��  ���        ���� � �����  �  s         ����  5 6           O^� � p     ����Pi  Y      �     ��  ���        ���� � �����  �  s         ����  7 8           Ve� � q     �����j  Xk   ��  �     ��  ���       ���� � �����  �  s         ����  9 :           ]l� � r     ���� l  �}   ��  �     ��  ���       ���� � �����  �  s         ����  ; <           ds� � s     �����m  �   ��  �     ��  ���       ���� � �����  �  s         ����  > ?           kz� � t     �����n  0�   ��  �     ��  ���       ����  �����  �  s         ����  @ A           r�� � u     ����Xp  x�   ��  �     ��  ���       ���� �����  �  s         ����  B C           y�� � v     �����q  ��   ��  �     ��  ���       ���� �����  �  s         ����  D E           ��� � w     ����(s  �   ��  �	     ��  ���       ���� �����  �  s         ����
  0 1           AH� � n     ����q  ��      ~      ��  ���        ���� � �����  �  t         ����
  2 3           HO� � o     ����tr  ��      ~     ��  ���        ���� � �����  �  t         ����
  4 5           OV� � p     �����s  ,�      ~     ��  ���        ���� � �����  �  t         ����
  6 7           V]� � q     ����Du  t�   ��  ~     ��  ���       ���� � �����  �  t         ����
  8 9           ]d� � r     �����v  �   ��  ~     ��  ���       ���� � �����  �  t         ����
  : ;           dk� � s     ����x     ��  ~     ��  ���       ���� � �����  �  t         ����
  = >           kr� � t     ����|y  L+   ��  ~     ��  ���       ����  �����  �  t         ����
  ? @           ry� � u     �����z  �=   ��  ~     ��  ���       ���� �����  �  t         ����
  A B           y�� � v     ����L|  �O   ��  ~     ��  ���       ���� �����  �  t         ����
  C D           ��� � w     �����}  $b   ��  ~	     ��  ���       ���� �����  �  t           ��  0 1           AT� � �     ����|o  L�             �     �        ���� � �����  �  u           ��  2 3           H[� � �     �����p  ��            �     �        ���� � �����  �  u           ��  4 5           Ob� � �     ����Lr  ��            �     �        ���� � �����  �  u         ! ��  6 7           Vi� � �     �����s  $�            �     �        ���� � �����  �  u         ! ��  8 9           ]p� � �     ����u  l�            �     �        ���� � �����  �  u         ! ��  : ;           dw� � �     �����v  �            �     �        ���� � �����  �  u         " ��  = >           k~� � �     �����w  �            �     �        ����  �����  �  u         " ��  ? @           r�� � �     ����Ty  D)            �     �        ���� �����  �  u         " ��  A B           y�� � �     �����z  �;            �     �        ���� �����  �  u         # ��  C D           ��� � �     ����$|  �M       	     �     �        ���� �����  �  u         ����  1 2           AZ� � n     �����u  ��      �      ��  ���        ���� � �����  �  v         ����  3 4           Ha� � o     ����$w  �      �     ��  ���        ���� � �����  �  v         ����  5 6           Oh� � p     �����x        �     ��  ���        ���� � �����  �  v         ����  7 8           Vo� � q     �����y  d1   ��  �     ��  ���       ���� � �����  �  v         ����  9 :           ]v� � r     ����\{  �C   ��  �     ��  ���       ���� � �����  �  v         ����  ; <           d}� � s     �����|  �U   ��  �     ��  ���       ���� � �����  �  v         ����  > ?           k�� � t     ����,~  <h   ��  �     ��  ���       ����  �����  �  v         ����  @ A           r�� � u     �����  �z   ��  �     ��  ���       ���� �����  �  v         ����  B C           y�� � v     ������  ̌   ��  �     ��  ���       ���� �����  �  v         ����  D E           ��� � w     ����d�  �   ��  �	     ��  ���       ���� �����  �  v         ����	  / 0           A@� � n     �����r  ��      $      ��  ���        ���� � �����  �  w         ����	  1 2           HG� � o     ����t  4�      $     ��  ���        ���� � �����  �  w         ����	  3 4           ON� � p     ����lu  |�      $     ��  ���        ���� � �����  �  w         ����	  5 6           VU� � q     �����v  �   ��  $     ��  ���       ���� � �����  �  w         ����	  7 8           ]\� � r     ����<x     ��  $     ��  ���       ���� � �����  �  w         ����	  9 :           dc� � s     �����y  T-   ��  $     ��  ���       ���� � �����  �  w         ����	  < =           kj� � t     ����{  �?   ��  $     ��  ���       ����  �����  �  w         ����	  > ?           rq� � u     ����t|  �Q   ��  $     ��  ���       ���� �����  �  w         ����	  @ A           yx� � v     �����}  ,d   ��  $     ��  ���       ���� �����  �  w         ����	  B C           �� � w     ����D  tv   ��  $	     ��  ���       ���� �����  �  w         ����  1 2           AX� � n     ����,t  <�      2      ��  ���        ���� � �����  �  x         ����  3 4           H_� � o     �����u  ��      2     ��  ���        ���� � �����  �  x         ����  5 6           Of� � p     �����v  �
      2     ��  ���        ���� � �����  �  x         ����  7 8           Vm� � q     ����dx     ��  2     ��  ���       ���� � �����  �  x         ����  9 :           ]t� � r     �����y  \/   ��  2     ��  ���       ���� � �����  �  x         ����  ; <           d{� � s     ����4{  �A   ��  2     ��  ���       ���� � �����  �  x         ����  > ?           k�� � t     �����|  �S   ��  2     ��  ���       ����  �����  �  x         ����  @ A           r�� � u     ����~  4f   ��  2     ��  ���       ���� �����  �  x         ����  B C           y�� � v     ����l  |x   ��  2     ��  ���       ���� �����  �  x         ����  D E           ��� � w     ����Ԁ  Ċ   ��  2	     ��  ���       ���� �����  �  x         ����   < =          �� � � n     z  �g  �C      !        ���        ���� � �����  �  y         ����   > ?          �� � o     �  i  V      !       ���        ���� � �����  �  y         ����   @ A          �� � p     �  |j  Lh      !       ���        ���� � �����  �  y         ����   C D          �� � q       �k  �z   ��  !       ���       ���� � �����  �  y         ����   E F          �� � r     5  Lm  ܌   ��  !       ���       ���� � �����  �  y         ����   G H          �� � s     d  �n  $�   ��  !       ���       ���� � �����  �  y         ����   I J          �� � t     �  p  l�   ��  !       ���       ����  �����  �  y         ����   K L          �%� � u     �  �q  ��   ��  !       ���       ���� �����  �  y         ����   N O          �+� � v     �  �r  ��   ��  !       ���       ���� �����  �  y         ����   P Q          �1� � w       Tt  D�   ��  !	       ���       ���� A  �  �  y         ����  ; <          �� � � n     ,  Te  D%      �        ���        ���� � �����  �  z         ����  = >          �� � o     [  �f  �7      �       ���        ���� � �����  �  z         ����  ? @          �� � p     �  $h  �I      �       ���        ���� � �����  �  z         ����  B C          �� � q     �  �i  \   ��  �       ���       ���� � �����  �  z         ����  D E          �� � r     �  �j  dn   ��  �       ���       ���� � �����  �  z         ����  F G          �� � s       \l  ��   ��  �       ���       ���� � �����  �  z         ����  H I          �� � t     E  �m  ��   ��  �       ���       ����  �����  �  z         ����  J K          �%� � u     s  ,o  <�   ��  �       ���       ���� �����  �  z         ����  M N          �+� � v     �  �p  ��   ��  �       ���       ���� �����  �  z         ����  O P          �1� � w     �  �q  ��   ��  �	       ���       ���� A  �  �  z         ����  : ;          �� � � n     9  �e  X*      �        ���        ���� � �����  �  {         ����  < =          �� � o     h   g  �<      �       ���        ���� � �����  �  {         ����  > ?          �� � p     �  �h  �N      �       ���        ���� � �����  �  {         ����  A B          �� � q     �  �i  0a   ��  �       ���       ���� � �����  �  {         ����  C D          �� � r     �  Xk  xs   ��  �       ���       ���� � �����  �  {         ����  E F          �� � s     #  �l  ��   ��  �       ���       ���� � �����  �  {         ����  G H          �� � t     R  (n  �   ��  �       ���       ����  �����  �  {         ����  I J          �%� � u     �  �o  P�   ��  �       ���       ���� �����  �  {         ����  L M          �+� � v     �  �p  ��   ��  �       ���       ���� �����  �  {         ����  N O          �1� � w     �  `r  ��   ��  �	       ���       ���� A  �  �  {         ����  : ;          �� � � n       \l  ��      a        ���        ���� � �����  �  |         ����  < =          �� � o     E  �m  ��      a       ���        ���� � �����  �  |         ����  > ?          �� � p     s  ,o  <�      a       ���        ���� � �����  �  |         ����  A B          �� � q     �  �p  ��   ��  a       ���       ���� � �����  �  |         ����  C D          �� � r     �  �q  ��   ��  a       ���       ���� � �����  �  |         ����  E F          �� � s        ds  �   ��  a       ���       ���� � �����  �  |         ����  G H          �� � t     /  �t  \�   ��  a       ���       ����  �����  �  |         ����  I J          �%� � u     ]  4v  �    ��  a       ���       ���� �����  �  |         ����  L M          �+� � v     �  �w  �   ��  a       ���       ���� �����  �  |         ����  N O          �1� � w     �  y  4%   ��  a	       ���       ���� A  �  �  |         ����  ; <          �� � � n     �  <i  X      -        ���        ���� � �����  �  }         ����  = >          �� � o     �  �j  Tj      -       ���        ���� � �����  �  }         ����  ? @          �� � p       l  �|      -       ���        ���� � �����  �  }         ����  B C          �� � q     :  tm  �   ��  -       ���       ���� � �����  �  }         ����  D E          �� � r     i  �n  ,�   ��  -       ���       ���� � �����  �  }         ����  F G          �� � s     �  Dp  t�   ��  -       ���       ���� � �����  �  }         ����  H I          �� � t     �  �q  ��   ��  -       ���       ����  �����  �  }         ����  J K          �%� � u     �  s  �   ��  -       ���       ���� �����  �  }         ����  M N          �+� � v     $  |t  L�   ��  -       ���       ���� �����  �  }         ����  O P          �1� � w     S  �u  ��   ��  -	       ���       ���� A  �  �  }         ����  = >          �� � � n     �  �j  \l      �        ���        ���� � �����  �  ~         ����  ? @          �� � o       4l  �~      �       ���        ���� � �����  �  ~         ����  A B          �� � p     ?  �m  �      �       ���        ���� � �����  �  ~         ����  D E          �� � q     n  o  4�   ��  �       ���       ���� � �����  �  ~         ����  F G          �� � r     �  lp  |�   ��  �       ���       ���� � �����  �  ~         ����  H I          �� � s     �  �q  ��   ��  �       ���       ���� � �����  �  ~         ����  J K          �� � t     �  <s  �   ��  �       ���       ����  �����  �  ~         ����  L M          �%� � u     )  �t  T�   ��  �       ���       ���� �����  �  ~         ����  O P          �+� � v     X  v  ��   ��  �       ���       ���� �����  �  ~         ����  Q R          �1� � w     �  tw  �   ��  �	       ���       ���� A  �  �  ~         ����  < =          �� � � n     J  �m  ��      �      �   �        ���� � �����  �           ����  > ?          �� � o     y  To  D�      �     �   �        ���� � �����  �           ����  @ A          �� � p     �  �p  ��      �     �   �        ���� � �����  �           ����  C D          �� � q     �  $r  ��   ��  �     �   �       ���� � �����  �           ����  E F          �� � r       �s  �   ��  �     �   �       ���� � �����  �           ����  G H          �� � s     4  �t  d�   ��  �     �   �       ���� � �����  �           ����  I J          �� � t     c  \v  �   ��  �     �   �       ����  �����  �           ����  K L          �%� � u     �  �w  �   ��  �     �   �       ���� �����  �           ����  N O          �+� � v     �  ,y  <'   ��  �     �   �       ���� �����  �           ����  P Q          �1� � w     �  �z  �9   ��  �	     �   �       ���� A  �  �           ����  < =           �� � � n     �����f  �4      �      �� ���        ���� � �����  �  �         ����  > ?           �� � o     �����g  �F      �     �� ���        ���� � �����  �  �         ����  @ A           �� � p     ����Pi  Y      �     �� ���        ���� � �����  �  �         ����  C D           �� � q     �����j  Xk   ��  �     �� ���       ���� � �����  �  �         ����  E F           �� � r     ���� l  �}   ��  �     �� ���       ���� � �����  �  �         ����  G H           �� � s     �����m  �   ��  �     �� ���       ���� � �����  �  �         ����  I J           �� � t     �����n  0�   ��  �     �� ���       ����  �����  �  �         ����  K L           �%� � u     ����Xp  x�   ��  �     �� ���       ���� �����  �  �         ����  N O           �+� � v     �����q  ��   ��  �     �� ���       ���� �����  �  �         ����  P Q           �1� � w     ����(s  �   ��  �	     �� ���       ���� �����  �  �         ����
  ; <           �� � � n     ����q  ��      B      �� ���        ���� � �����  �  �         ����
  = >           �� � o     ����tr  ��      B     �� ���        ���� � �����  �  �         ����
  ? @           �� � p     �����s  ,�      B     �� ���        ���� � �����  �  �         ����
  B C           �� � q     ����Du  t�   ��  B     �� ���       ���� � �����  �  �         ����
  D E           �� � r     �����v  �   ��  B     �� ���       ���� � �����  �  �         ����
  F G           �� � s     ����x     ��  B     �� ���       ���� � �����  �  �         ����
  H I           �� � t     ����|y  L+   ��  B     �� ���       ����  �����  �  �         ����
  J K           �%� � u     �����z  �=   ��  B     �� ���       ���� �����  �  �         ����
  M N           �+� � v     ����L|  �O   ��  B     �� ���       ���� �����  �  �         ����
  O P           �1� � w     �����}  $b   ��  B	     �� ���       ���� �����  �  �           ��  = >           �� � � �     ����|o  L�       �       �    �        ���� � �����  �  �           ��  ? @           �� � �     �����p  ��       �      �    �        ���� � �����  �  �           ��  A B           �� � �     ����Lr  ��       �      �    �        ���� � �����  �  �         ! ��  D E           �� � �     �����s  $�       �      �    �        ���� � �����  �  �         ! ��  F G           �� � �     ����u  l�       �      �    �        ���� � �����  �  �         ! ��  H I           �� � �     �����v  �       �      �    �        ���� � �����  �  �         " ��  J K           �� � �     �����w  �       �      �    �        ����  �����  �  �         " ��  L M           �%� � �     ����Ty  D)       �      �    �        ���� �����  �  �         " ��  O P           �+� � �     �����z  �;       �      �    �        ���� �����  �  �         # ��  Q R           1� � �     ����$|  �M       � 	     �    �        ���� �����  �  �         ����  = >           �� � � n     �����u  ��      P      �� ���        ���� � �����  �  �         ����  ? @           �� � o     ����$w  �      P     �� ���        ���� � �����  �  �         ����  A B           �� � p     �����x        P     �� ���        ���� � �����  �  �         ����  D E           �� � q     �����y  d1   ��  P     �� ���       ���� � �����  �  �         ����  F G           �� � r     ����\{  �C   ��  P     �� ���       ���� � �����  �  �         ����  H I           �� � s     �����|  �U   ��  P     �� ���       ���� � �����  �  �         ����  J K           �� � t     ����,~  <h   ��  P     �� ���       ����  �����  �  �         ����  L M           �%� � u     �����  �z   ��  P     �� ���       ���� �����  �  �         ����  O P           �+� � v     ������  ̌   ��  P     �� ���       ���� �����  �  �         ����  Q R           1� � w     ����d�  �   ��  P	     �� ���       ���� �����  �  �         ����	  : ;           �� � � n     �����r  ��      �      �� ���        ���� � �����  �  �         ����	  < =           �� � o     ����t  4�      �     �� ���        ���� � �����  �  �         ����	  > ?           �� � p     ����lu  |�      �     �� ���        ���� � �����  �  �         ����	  A B           �� � q     �����v  �   ��  �     �� ���       ���� � �����  �  �         ����	  C D           �� � r     ����<x     ��  �     �� ���       ���� � �����  �  �         ����	  E F           �� � s     �����y  T-   ��  �     �� ���       ���� � �����  �  �         ����	  G H           �� � t     ����{  �?   ��  �     �� ���       ����  �����  �  �         ����	  I J           �%� � u     ����t|  �Q   ��  �     �� ���       ���� �����  �  �         ����	  L M           �+� � v     �����}  ,d   ��  �     �� ���       ���� �����  �  �         ����	  N O           �1� � w     ����D  tv   ��  �	     �� ���       ���� �����  �  �         ����  = >           �� � � n     ����,t  <�      �      �� ���        ���� � �����  �  �         ����  ? @           �� � o     �����u  ��      �     �� ���        ���� � �����  �  �         ����  A B           �� � p     �����v  �
      �     �� ���        ���� � �����  �  �         ����  D E           �� � q     ����dx     ��  �     �� ���       ���� � �����  �  �         ����  F G           �� � r     �����y  \/   ��  �     �� ���       ���� � �����  �  �         ����  H I           �� � s     ����4{  �A   ��  �     �� ���       ���� � �����  �  �         ����  J K           �� � t     �����|  �S   ��  �     �� ���       ����  �����  �  �         ����  L M           �%� � u     ����~  4f   ��  �     �� ���       ���� �����  �  �         ����  O P           �+� � v     ����l  |x   ��  �     �� ���       ���� �����  �  �         ����  Q R           1� � w     ����Ԁ  Ċ   ��  �	     �� ���       ���� �����  �  �         ����   / 0          � � �� n     z  �g  �C      5        ���        ���� � �����  �  �         ����   1 2          � � �� o     �  i  V      5       ���        ���� � �����  �  �         ����   3 4          � �� p     �  |j  Lh      5       ���        ���� � �����  �  �         ����   5 6          � 	�� q       �k  �z   ��  5       ���       ���� � �����  �  �         ����   7 8          � �� r     5  Lm  ܌   ��  5       ���       ���� � �����  �  �         ����   9 :          � �� s     d  �n  $�   ��  5       ���       ���� � �����  �  �         ����   < =          � �� t     �  p  l�   ��  5       ���       ����  �����  �  �         ����   > ?          � !�� u     �  �q  ��   ��  5       ���       ���� �����  �  �         ����   @ A          � '�� v     �  �r  ��   ��  5       ���       ���� �����  �  �         ����   B C          � -�� w       Tt  D�   ��  5	       ���       ���� A  �  �  �         ����  . /          � � �� n     ,  Te  D%              ���        ���� � �����  �  �         ����  0 1          � � �� o     [  �f  �7             ���        ���� � �����  �  �         ����  2 3          � � �� p     �  $h  �I             ���        ���� � �����  �  �         ����  4 5          � �� q     �  �i  \   ��         ���       ���� � �����  �  �         ����  6 7          � �� r     �  �j  dn   ��         ���       ���� � �����  �  �         ����  8 9          � �� s       \l  ��   ��         ���       ���� � �����  �  �         ����  ; <          � �� t     E  �m  ��   ��         ���       ����  �����  �  �         ����  = >          � �� u     s  ,o  <�   ��         ���       ���� �����  �  �         ����  ? @          � �� v     �  �p  ��   ��         ���       ���� �����  �  �         ����  A B          � %�� w     �  �q  ��   ��  	       ���       ���� A  �  �  �         ����  . /          � � �� n     9  �e  X*      �        ���        ���� � �����  �  �         ����  0 1          � � �� o     h   g  �<      �       ���        ���� � �����  �  �         ����  2 3          � � �� p     �  �h  �N      �       ���        ���� � �����  �  �         ����  4 5          � � �� q     �  �i  0a   ��  �       ���       ���� � �����  �  �         ����  6 7          � � �� r     �  Xk  xs   ��  �       ���       ���� � �����  �  �         ����  8 9          �  �� s     #  �l  ��   ��  �       ���       ���� � �����  �  �         ����  ; <          � �� t     R  (n  �   ��  �       ���       ����  �����  �  �         ����  = >          � �� u     �  �o  P�   ��  �       ���       ���� �����  �  �         ����  ? @          � �� v     �  �p  ��   ��  �       ���       ���� �����  �  �         ����  A B          � �� w     �  `r  ��   ��  �	       ���       ���� A  �  �  �         ����  . /          � � �� n       \l  ��      r        ���        ���� � �����  �  �         ����  0 1          � � �� o     E  �m  ��      r       ���        ���� � �����  �  �         ����  2 3          � � �� p     s  ,o  <�      r       ���        ���� � �����  �  �         ����  4 5          � � �� q     �  �p  ��   ��  r       ���       ���� � �����  �  �         ����  6 7          � � �� r     �  �q  ��   ��  r       ���       ���� � �����  �  �         ����  8 9          � � �� s        ds  �   ��  r       ���       ���� � �����  �  �         ����  ; <          � �� t     /  �t  \�   ��  r       ���       ����  �����  �  �         ����  = >          � �� u     ]  4v  �    ��  r       ���       ���� �����  �  �         ����  ? @          � �� v     �  �w  �   ��  r       ���       ���� �����  �  �         ����  A B          � �� w     �  y  4%   ��  r	       ���       ���� A  �  �  �         ����  . /          � � �� n     �  <i  X      >        ���        ���� � �����  �  �         ����  0 1          � � �� o     �  �j  Tj      >       ���        ���� � �����  �  �         ����  2 3          � � �� p       l  �|      >       ���        ���� � �����  �  �         ����  4 5          � � �� q     :  tm  �   ��  >       ���       ���� � �����  �  �         ����  6 7          � �� r     i  �n  ,�   ��  >       ���       ���� � �����  �  �         ����  8 9          � �� s     �  Dp  t�   ��  >       ���       ���� � �����  �  �         ����  ; <          � �� t     �  �q  ��   ��  >       ���       ����  �����  �  �         ����  = >          � �� u     �  s  �   ��  >       ���       ���� �����  �  �         ����  ? @          � �� v     $  |t  L�   ��  >       ���       ���� �����  �  �         ����  A B          �  �� w     S  �u  ��   ��  >	       ���       ���� A  �  �  �         ����  / 0          � �� n     �  �j  \l      �        ���        ���� � �����  �  �         ����  1 2          � 
�� o       4l  �~      �       ���        ���� � �����  �  �         ����  3 4          � �� p     ?  �m  �      �       ���        ���� � �����  �  �         ����  5 6          � �� q     n  o  4�   ��  �       ���       ���� � �����  �  �         ����  7 8          � �� r     �  lp  |�   ��  �       ���       ���� � �����  �  �         ����  9 :          � "�� s     �  �q  ��   ��  �       ���       ���� � �����  �  �         ����  < =          � (�� t     �  <s  �   ��  �       ���       ����  �����  �  �         ����  > ?          � .�� u     )  �t  T�   ��  �       ���       ���� �����  �  �         ����  @ A          � 4�� v     X  v  ��   ��  �       ���       ���� �����  �  �         ����  B C          � :�� w     �  tw  �   ��  �	       ���       ���� A  �  �  �         ����  / 0          � � �� n     J  �m  ��      �      �   �        ���� � �����  �  �         ����  1 2          � �� o     y  To  D�      �     �   �        ���� � �����  �  �         ����  3 4          � �� p     �  �p  ��      �     �   �        ���� � �����  �  �         ����  5 6          � �� q     �  $r  ��   ��  �     �   �       ���� � �����  �  �         ����  7 8          � �� r       �s  �   ��  �     �   �       ���� � �����  �  �         ����  9 :          � �� s     4  �t  d�   ��  �     �   �       ���� � �����  �  �         ����  < =          �  �� t     c  \v  �   ��  �     �   �       ����  �����  �  �         ����  > ?          � &�� u     �  �w  �   ��  �     �   �       ���� �����  �  �         ����  @ A          � ,�� v     �  ,y  <'   ��  �     �   �       ���� �����  �  �         ����  B C          � 2�� w     �  �z  �9   ��  �	     �   �       ���� A  �  �  �         ����  / 0           � � �� n     �����f  �4      �      �� ���        ���� � �����  �  �         ����  1 2           � �� o     �����g  �F      �     �� ���        ���� � �����  �  �         ����  3 4           � �� p     ����Pi  Y      �     �� ���        ���� � �����  �  �         ����  5 6           � �� q     �����j  Xk   ��  �     �� ���       ���� � �����  �  �         ����  7 8           � �� r     ���� l  �}   ��  �     �� ���       ���� � �����  �  �         ����  9 :           � �� s     �����m  �   ��  �     �� ���       ���� � �����  �  �         ����  < =           � #�� t     �����n  0�   ��  �     �� ���       ����  �����  �  �         ����  > ?           � )�� u     ����Xp  x�   ��  �     �� ���       ���� �����  �  �         ����  @ A           � /�� v     �����q  ��   ��  �     �� ���       ���� �����  �  �         ����  B C           � 5�� w     ����(s  �   ��  �	     �� ���       ���� �����  �  �         ����
  . /           � � �� n     ����q  ��      Q      �� ���        ���� � �����  �  �         ����
  0 1           � � �� o     ����tr  ��      Q     �� ���        ���� � �����  �  �         ����
  2 3           � � �� p     �����s  ,�      Q     �� ���        ���� � �����  �  �         ����
  4 5           � �� q     ����Du  t�   ��  Q     �� ���       ���� � �����  �  �         ����
  6 7           � 
�� r     �����v  �   ��  Q     �� ���       ���� � �����  �  �         ����
  8 9           � �� s     ����x     ��  Q     �� ���       ���� � �����  �  �         ����
  ; <           � �� t     ����|y  L+   ��  Q     �� ���       ����  �����  �  �         ����
  = >           � �� u     �����z  �=   ��  Q     �� ���       ���� �����  �  �         ����
  ? @           � "�� v     ����L|  �O   ��  Q     �� ���       ���� �����  �  �         ����
  A B           � (�� w     �����}  $b   ��  Q	     �� ���       ���� �����  �  �           ��  / 0           � 	�� �     ����|o  L�       �       �    �        ���� � �����  �  �           ��  1 2           � �� �     �����p  ��       �      �    �        ���� � �����  �  �           ��  3 4           � �� �     ����Lr  ��       �      �    �        ���� � �����  �  �         ! ��  5 6           � �� �     �����s  $�       �      �    �        ���� � �����  �  �         ! ��  7 8           � !�� �     ����u  l�       �      �    �        ���� � �����  �  �         ! ��  9 :           � '�� �     �����v  �       �      �    �        ���� � �����  �  �         " ��  < =           � -�� �     �����w  �       �      �    �        ����  �����  �  �         " ��  > ?           � 3�� �     ����Ty  D)       �      �    �        ���� �����  �  �         " ��  @ A           � 9�� �     �����z  �;       �      �    �        ���� �����  �  �         # ��  B C           � ?�� �     ����$|  �M       � 	     �    �        ���� �����  �  �         ����  / 0           � �� n     �����u  ��      _      �� ���        ���� � �����  �  �         ����  1 2           � �� o     ����$w  �      _     �� ���        ���� � �����  �  �         ����  3 4           � �� p     �����x        _     �� ���        ���� � �����  �  �         ����  5 6           � !�� q     �����y  d1   ��  _     �� ���       ���� � �����  �  �         ����  7 8           � '�� r     ����\{  �C   ��  _     �� ���       ���� � �����  �  �         ����  9 :           � -�� s     �����|  �U   ��  _     �� ���       ���� � �����  �  �         ����  < =           � 3�� t     ����,~  <h   ��  _     �� ���       ����  �����  �  �         ����  > ?           � 9�� u     �����  �z   ��  _     �� ���       ���� �����  �  �         ����  @ A           � ?�� v     ������  ̌   ��  _     �� ���       ���� �����  �  �         ����  B C           � E � w     ����d�  �   ��  _	     �� ���       ���� �����  �  �         ����	  . /           � � �� n     �����r  ��      �      �� ���        ���� � �����  �  �         ����	  0 1           � � �� o     ����t  4�      �     �� ���        ���� � �����  �  �         ����	  2 3           � � �� p     ����lu  |�      �     �� ���        ���� � �����  �  �         ����	  4 5           � � �� q     �����v  �   ��  �     �� ���       ���� � �����  �  �         ����	  6 7           � � �� r     ����<x     ��  �     �� ���       ���� � �����  �  �         ����	  8 9           � �� s     �����y  T-   ��  �     �� ���       ���� � �����  �  �         ����	  ; <           � 	�� t     ����{  �?   ��  �     �� ���       ����  �����  �  �         ����	  = >           � �� u     ����t|  �Q   ��  �     �� ���       ���� �����  �  �         ����	  ? @           � �� v     �����}  ,d   ��  �     �� ���       ���� �����  �  �         ����	  A B           � �� w     ����D  tv   ��  �	     �� ���       ���� �����  �  �         ����  / 0           � �� n     ����,t  <�            �� ���        ���� � �����  �  �         ����  1 2           � �� o     �����u  ��           �� ���        ���� � �����  �  �         ����  3 4           � �� p     �����v  �
           �� ���        ���� � �����  �  �         ����  5 6           � �� q     ����dx     ��       �� ���       ���� � �����  �  �         ����  7 8           � $�� r     �����y  \/   ��       �� ���       ���� � �����  �  �         ����  9 :           � *�� s     ����4{  �A   ��       �� ���       ���� � �����  �  �         ����  < =           � 0�� t     �����|  �S   ��       �� ���       ����  �����  �  �         ����  > ?           � 6�� u     ����~  4f   ��       �� ���       ���� �����  �  �         ����  @ A           � <�� v     ����l  |x   ��       �� ���       ���� �����  �  �         ����  B C           � B�� w     ����Ԁ  Ċ   ��  	     �� ���       ���� �����  �  �         ����   . /          ]� ]� n     z  �g  �C      I        ���        ���� � �����  �  �         ����   0 1          d� d� o     �  i  V      I       ���        ���� � �����  �  �         ����   2 3          k� k� p     �  |j  Lh      I       ���        ���� � �����  �  �         ����   4 5          r� r� q       �k  �z   ��  I       ���       ���� � �����  �  �         ����   6 7          y� y� r     5  Lm  ܌   ��  I       ���       ���� � �����  �  �         ����   8 9          �� �� s     d  �n  $�   ��  I       ���       ���� � �����  �  �         ����   ; <          �� �� t     �  p  l�   ��  I       ���       ����  �����  �  �         ����   = >          �� �� u     �  �q  ��   ��  I       ���       ���� �����  �  �         ����   ? @          �� �� v     �  �r  ��   ��  I       ���       ���� �����  �  �         ����   A B          �� �� w       Tt  D�   ��  I	       ���       ���� A  �  �  �         ����  - .          U� U� n     ,  Te  D%              ���        ���� � �����  �  �         ����  / 0          \� \� o     [  �f  �7             ���        ���� � �����  �  �         ����  1 2          c� c� p     �  $h  �I             ���        ���� � �����  �  �         ����  3 4          j� j� q     �  �i  \   ��         ���       ���� � �����  �  �         ����  5 6          q� q� r     �  �j  dn   ��         ���       ���� � �����  �  �         ����  7 8          x� x� s       \l  ��   ��         ���       ���� � �����  �  �         ����  : ;          � � t     E  �m  ��   ��         ���       ����  �����  �  �         ����  < =          �� �� u     s  ,o  <�   ��         ���       ���� �����  �  �         ����  > ?          �� �� v     �  �p  ��   ��         ���       ���� �����  �  �         ����  @ A          �� �� w     �  �q  ��   ��  	       ���       ���� A  �  �  �         ����  - .          H� H� n     9  �e  X*      �        ���        ���� � �����  �  �         ����  / 0          O� O� o     h   g  �<      �       ���        ���� � �����  �  �         ����  1 2          V� V� p     �  �h  �N      �       ���        ���� � �����  �  �         ����  3 4          ]� ]� q     �  �i  0a   ��  �       ���       ���� � �����  �  �         ����  5 6          d� d� r     �  Xk  xs   ��  �       ���       ���� � �����  �  �         ����  7 8          k� k� s     #  �l  ��   ��  �       ���       ���� � �����  �  �         ����  : ;          r� r� t     R  (n  �   ��  �       ���       ����  �����  �  �         ����  < =          y� y� u     �  �o  P�   ��  �       ���       ���� �����  �  �         ����  > ?          �� �� v     �  �p  ��   ��  �       ���       ���� �����  �  �         ����  @ A          �� �� w     �  `r  ��   ��  �	       ���       ���� A  �  �  �         ����  - .          C� C� n       \l  ��      �        ���        ���� � �����  �  �         ����  / 0          J� J� o     E  �m  ��      �       ���        ���� � �����  �  �         ����  1 2          Q� Q� p     s  ,o  <�      �       ���        ���� � �����  �  �         ����  3 4          X� X� q     �  �p  ��   ��  �       ���       ���� � �����  �  �         ����  5 6          _� _� r     �  �q  ��   ��  �       ���       ���� � �����  �  �         ����  7 8          f� f� s        ds  �   ��  �       ���       ���� � �����  �  �         ����  : ;          m� m� t     /  �t  \�   ��  �       ���       ����  �����  �  �         ����  < =          t� t� u     ]  4v  �    ��  �       ���       ���� �����  �  �         ����  > ?          {� {� v     �  �w  �   ��  �       ���       ���� �����  �  �         ����  @ A          �� �� w     �  y  4%   ��  �	       ���       ���� A  �  �  �         ����  - .          P� P� n     �  <i  X      O        ���        ���� � �����  �  �         ����  / 0          W� W� o     �  �j  Tj      O       ���        ���� � �����  �  �         ����  1 2          ^� ^� p       l  �|      O       ���        ���� � �����  �  �         ����  3 4          e� e� q     :  tm  �   ��  O       ���       ���� � �����  �  �         ����  5 6          l� l� r     i  �n  ,�   ��  O       ���       ���� � �����  �  �         ����  7 8          s� s� s     �  Dp  t�   ��  O       ���       ���� � �����  �  �         ����  : ;          z� z� t     �  �q  ��   ��  O       ���       ����  �����  �  �         ����  < =          �� �� u     �  s  �   ��  O       ���       ���� �����  �  �         ����  > ?          �� �� v     $  |t  L�   ��  O       ���       ���� �����  �  �         ����  @ A          �� �� w     S  �u  ��   ��  O	       ���       ���� A  �  �  �         ����  . /          j� j� n     �  �j  \l      �        ���        ���� � �����  �  �         ����  0 1          q� q� o       4l  �~      �       ���        ���� � �����  �  �         ����  2 3          x� x� p     ?  �m  �      �       ���        ���� � �����  �  �         ����  4 5          � � q     n  o  4�   ��  �       ���       ���� � �����  �  �         ����  6 7          �� �� r     �  lp  |�   ��  �       ���       ���� � �����  �  �         ����  8 9          �� �� s     �  �q  ��   ��  �       ���       ���� � �����  �  �         ����  ; <          �� �� t     �  <s  �   ��  �       ���       ����  �����  �  �         ����  = >          �� �� u     )  �t  T�   ��  �       ���       ���� �����  �  �         ����  ? @          �� �� v     X  v  ��   ��  �       ���       ���� �����  �  �         ����  A B          �� �� w     �  tw  �   ��  �	       ���       ���� A  �  �  �         ����  . /          b� b� n     J  �m  ��      �      �   �        ���� � �����  �  �         ����  0 1          i� i� o     y  To  D�      �     �   �        ���� � �����  �  �         ����  2 3          p� p� p     �  �p  ��      �     �   �        ���� � �����  �  �         ����  4 5          w� w� q     �  $r  ��   ��  �     �   �       ���� � �����  �  �         ����  6 7          ~� ~� r       �s  �   ��  �     �   �       ���� � �����  �  �         ����  8 9          �� �� s     4  �t  d�   ��  �     �   �       ���� � �����  �  �         ����  ; <          �� �� t     c  \v  �   ��  �     �   �       ����  �����  �  �         ����  = >          �� �� u     �  �w  �   ��  �     �   �       ���� �����  �  �         ����  ? @          �� �� v     �  ,y  <'   ��  �     �   �       ���� �����  �  �         ����  A B          �� �� w     �  �z  �9   ��  �	     �   �       ���� A  �  �  �         ����  . /           e� e� n     �����f  �4      �      �� ���        ���� � �����  �  �         ����  0 1           l� l� o     �����g  �F      �     �� ���        ���� � �����  �  �         ����  2 3           s� s� p     ����Pi  Y      �     �� ���        ���� � �����  �  �         ����  4 5           z� z� q     �����j  Xk   ��  �     �� ���       ���� � �����  �  �         ����  6 7           �� �� r     ���� l  �}   ��  �     �� ���       ���� � �����  �  �         ����  8 9           �� �� s     �����m  �   ��  �     �� ���       ���� � �����  �  �         ����  ; <           �� �� t     �����n  0�   ��  �     �� ���       ����  �����  �  �         ����  = >           �� �� u     ����Xp  x�   ��  �     �� ���       ���� �����  �  �         ����  ? @           �� �� v     �����q  ��   ��  �     �� ���       ���� �����  �  �         ����  A B           �� �� w     ����(s  �   ��  �	     �� ���       ���� �����  �  �         ����
  - .           X� X� n     ����q  ��      `      �� ���        ���� � �����  �  �         ����
  / 0           _� _� o     ����tr  ��      `     �� ���        ���� � �����  �  �         ����
  1 2           f� f� p     �����s  ,�      `     �� ���        ���� � �����  �  �         ����
  3 4           m� m� q     ����Du  t�   ��  `     �� ���       ���� � �����  �  �         ����
  5 6           t� t� r     �����v  �   ��  `     �� ���       ���� � �����  �  �         ����
  7 8           {� {� s     ����x     ��  `     �� ���       ���� � �����  �  �         ����
  : ;           �� �� t     ����|y  L+   ��  `     �� ���       ����  �����  �  �         ����
  < =           �� �� u     �����z  �=   ��  `     �� ���       ���� �����  �  �         ����
  > ?           �� �� v     ����L|  �O   ��  `     �� ���       ���� �����  �  �         ����
  @ A           �� �� w     �����}  $b   ��  `	     �� ���       ���� �����  �  �           ��  . /           o� o� �     ����|o  L�       �       �    �        ���� � �����  �  �           ��  0 1           v� v� �     �����p  ��       �      �    �        ���� � �����  �  �           ��  2 3           }� }� �     ����Lr  ��       �      �    �        ���� � �����  �  �         ! ��  4 5           �� �� �     �����s  $�       �      �    �        ���� � �����  �  �         ! ��  6 7           �� �� �     ����u  l�       �      �    �        ���� � �����  �  �         ! ��  8 9           �� �� �     �����v  �       �      �    �        ���� � �����  �  �         " ��  ; <           �� �� �     �����w  �       �      �    �        ����  �����  �  �         " ��  = >           �� �� �     ����Ty  D)       �      �    �        ���� �����  �  �         " ��  ? @           �� �� �     �����z  �;       �      �    �        ���� �����  �  �         # ��  A B           �� �� �     ����$|  �M       � 	     �    �        ���� �����  �  �         ����  . /           u� u� n     �����u  ��      n      �� ���        ���� � �����  �  �         ����  0 1           |� |� o     ����$w  �      n     �� ���        ���� � �����  �  �         ����  2 3           �� �� p     �����x        n     �� ���        ���� � �����  �  �         ����  4 5           �� �� q     �����y  d1   ��  n     �� ���       ���� � �����  �  �         ����  6 7           �� �� r     ����\{  �C   ��  n     �� ���       ���� � �����  �  �         ����  8 9           �� �� s     �����|  �U   ��  n     �� ���       ���� � �����  �  �         ����  ; <           �� �� t     ����,~  <h   ��  n     �� ���       ����  �����  �  �         ����  = >           �� �� u     �����  �z   ��  n     �� ���       ���� �����  �  �         ����  ? @           �� �� v     ������  ̌   ��  n     �� ���       ���� �����  �  �         ����  A B           �� �� w     ����d�  �   ��  n	     �� ���       ���� �����  �  �         ����	  - .           K� K� n     �����r  ��            �� ���        ���� � �����  �  �         ����	  / 0           R� R� o     ����t  4�           �� ���        ���� � �����  �  �         ����	  1 2           Y� Y� p     ����lu  |�           �� ���        ���� � �����  �  �         ����	  3 4           `� `� q     �����v  �   ��       �� ���       ���� � �����  �  �         ����	  5 6           g� g� r     ����<x     ��       �� ���       ���� � �����  �  �         ����	  7 8           n� n� s     �����y  T-   ��       �� ���       ���� � �����  �  �         ����	  : ;           u� u� t     ����{  �?   ��       �� ���       ����  �����  �  �         ����	  < =           |� |� u     ����t|  �Q   ��       �� ���       ���� �����  �  �         ����	  > ?           �� �� v     �����}  ,d   ��       �� ���       ���� �����  �  �         ����	  @ A           �� �� w     ����D  tv   ��  	     �� ���       ���� �����  �  �         ����  . /           r� r� n     ����,t  <�            �� ���        ���� � �����  �  �         ����  0 1           y� y� o     �����u  ��           �� ���        ���� � �����  �  �         ����  2 3           �� �� p     �����v  �
           �� ���        ���� � �����  �  �         ����  4 5           �� �� q     ����dx     ��       �� ���       ���� � �����  �  �         ����  6 7           �� �� r     �����y  \/   ��       �� ���       ���� � �����  �  �         ����  8 9           �� �� s     ����4{  �A   ��       �� ���       ���� � �����  �  �         ����  ; <           �� �� t     �����|  �S   ��       �� ���       ����  �����  �  �         ����  = >           �� �� u     ����~  4f   ��       �� ���       ���� �����  �  �         ����  ? @           �� �� v     ����l  |x   ��       �� ���       ���� �����  �  �         ����  A B           �� �� w     ����Ԁ  Ċ   ��  	     �� ���       ���� �����  �  �         ����   # $          � � �� n     z  �g  �C      ]        ���        ���� � �����  �  �         ����   % &          � � �� o     �  i  V      ]       ���        ���� � �����  �  �         ����   ' (          � � �� p     �  |j  Lh      ]       ���        ���� � �����  �  �         ����   ) *          � � �� q       �k  �z   ��  ]       ���       ���� � �����  �  �         ����   + ,          � �� r     5  Lm  ܌   ��  ]       ���       ���� � �����  �  �         ����   - .          � 
�� s     d  �n  $�   ��  ]       ���       ���� � �����  �  �         ����   / 0          � �� t     �  p  l�   ��  ]       ���       ����  �����  �  �         ����   1 2          � �� u     �  �q  ��   ��  ]       ���       ���� �����  �  �         ����   3 4          � �� v     �  �r  ��   ��  ]       ���       ���� �����  �  �         ����   5 6          � "�� w       Tt  D�   ��  ]	       ���       ���� A  �  �  �         ����  " #          � � �� n     ,  Te  D%      .        ���        ���� � �����  �  �         ����  $ %          � � �� o     [  �f  �7      .       ���        ���� � �����  �  �         ����  & '          � � �� p     �  $h  �I      .       ���        ���� � �����  �  �         ����  ( )          �  �� q     �  �i  \   ��  .       ���       ���� � �����  �  �         ����  * +          � �� r     �  �j  dn   ��  .       ���       ���� � �����  �  �         ����  , -          � �� s       \l  ��   ��  .       ���       ���� � �����  �  �         ����  . /          � �� t     E  �m  ��   ��  .       ���       ����  �����  �  �         ����  0 1          � �� u     s  ,o  <�   ��  .       ���       ���� �����  �  �         ����  2 3          � �� v     �  �p  ��   ��  .       ���       ���� �����  �  �         ����  4 5          � $�� w     �  �q  ��   ��  .	       ���       ���� A  �  �  �         ����  " #          � � �� n     9  �e  X*      �        ���        ���� � �����  �  �         ����  $ %          � � �� o     h   g  �<      �       ���        ���� � �����  �  �         ����  & '          � � �� p     �  �h  �N      �       ���        ���� � �����  �  �         ����  ( )          � � �� q     �  �i  0a   ��  �       ���       ���� � �����  �  �         ����  * +          � � �� r     �  Xk  xs   ��  �       ���       ���� � �����  �  �         ����  , -          � �� s     #  �l  ��   ��  �       ���       ���� � �����  �  �         ����  . /          � �� t     R  (n  �   ��  �       ���       ����  �����  �  �         ����  0 1          � �� u     �  �o  P�   ��  �       ���       ���� �����  �  �         ����  2 3          � �� v     �  �p  ��   ��  �       ���       ���� �����  �  �         ����  4 5          � �� w     �  `r  ��   ��  �	       ���       ���� A  �  �  �         ����  " #          � � �} n       \l  ��      �        ���        ���� � �����  �  �         ����  $ %          � � �� o     E  �m  ��      �       ���        ���� � �����  �  �         ����  & '          � � �� p     s  ,o  <�      �       ���        ���� � �����  �  �         ����  ( )          � � �� q     �  �p  ��   ��  �       ���       ���� � �����  �  �         ����  * +          � � �� r     �  �q  ��   ��  �       ���       ���� � �����  �  �         ����  , -          � � �� s        ds  �   ��  �       ���       ���� � �����  �  �         ����  . /          � �� t     /  �t  \�   ��  �       ���       ����  �����  �  �         ����  0 1          � 
�� u     ]  4v  �    ��  �       ���       ���� �����  �  �         ����  2 3          � �� v     �  �w  �   ��  �       ���       ���� �����  �  �         ����  4 5          � �� w     �  y  4%   ��  �	       ���       ���� A  �  �  �         ����  " #          � � �� n     �  <i  X      `        ���        ���� � �����  �  �         ����  $ %          � � �� o     �  �j  Tj      `       ���        ���� � �����  �  �         ����  & '          � � �� p       l  �|      `       ���        ���� � �����  �  �         ����  ( )          � �� q     :  tm  �   ��  `       ���       ���� � �����  �  �         ����  * +          � 
�� r     i  �n  ,�   ��  `       ���       ���� � �����  �  �         ����  , -          � �� s     �  Dp  t�   ��  `       ���       ���� � �����  �  �         ����  . /          � �� t     �  �q  ��   ��  `       ���       ����  �����  �  �         ����  0 1          � �� u     �  s  �   ��  `       ���       ���� �����  �  �         ����  2 3          � "�� v     $  |t  L�   ��  `       ���       ���� �����  �  �         ����  4 5          � (�� w     S  �u  ��   ��  `	       ���       ���� A  �  �  �         ����  # $          � � �� n     �  �j  \l      �        ���        ���� � �����  �  �         ����  % &          � �� o       4l  �~      �       ���        ���� � �����  �  �         ����  ' (          � �� p     ?  �m  �      �       ���        ���� � �����  �  �         ����  ) *          � �� q     n  o  4�   ��  �       ���       ���� � �����  �  �         ����  + ,          � �� r     �  lp  |�   ��  �       ���       ���� � �����  �  �         ����  - .          � �� s     �  �q  ��   ��  �       ���       ���� � �����  �  �         ����  / 0          � �� t     �  <s  �   ��  �       ���       ����  �����  �  �         ����  1 2          � %�� u     )  �t  T�   ��  �       ���       ���� �����  �  �         ����  3 4          � +�� v     X  v  ��   ��  �       ���       ���� �����  �  �         ����  5 6          � 1�� w     �  tw  �   ��  �	       ���       ���� A  �  �  �         ����  $ %          � � �� n     J  �m  ��      �      �   �        ���� � �����  �  �         ����  & '          � � �� o     y  To  D�      �     �   �        ���� � �����  �  �         ����  ( )          � � �� p     �  �p  ��      �     �   �        ���� � �����  �  �         ����  * +          � � �� q     �  $r  ��   ��  �     �   �       ���� � �����  �  �         ����  , -          � � �� r       �s  �   ��  �     �   �       ���� � �����  �  �         ����  . /          � � �� s     4  �t  d�   ��  �     �   �       ���� � �����  �  �         ����  0 1          � �� t     c  \v  �   ��  �     �   �       ����  �����  �  �         ����  2 3          � 	�� u     �  �w  �   ��  �     �   �       ���� �����  �  �         ����  4 5          � �� v     �  ,y  <'   ��  �     �   �       ���� �����  �  �         ����  6 7          � �� w     �  �z  �9   ��  �	     �   �       ���� A  �  �  �         ����  # $           � � �� n     �����f  �4      �      �� ���        ���� � �����  �  �         ����  % &           � � �� o     �����g  �F      �     �� ���        ���� � �����  �  �         ����  ' (           � � �� p     ����Pi  Y      �     �� ���        ���� � �����  �  �         ����  ) *           �  �� q     �����j  Xk   ��  �     �� ���       ���� � �����  �  �         ����  + ,           � �� r     ���� l  �}   ��  �     �� ���       ���� � �����  �  �         ����  - .           � �� s     �����m  �   ��  �     �� ���       ���� � �����  �  �         ����  / 0           � �� t     �����n  0�   ��  �     �� ���       ����  �����  �  �         ����  1 2           � �� u     ����Xp  x�   ��  �     �� ���       ���� �����  �  �         ����  3 4           � �� v     �����q  ��   ��  �     �� ���       ���� �����  �  �         ����  5 6           � $�� w     ����(s  �   ��  �	     �� ���       ���� �����  �  �         ����
  # $           � � �� n     ����q  ��      o      �� ���        ���� � �����  �  �         ����
  % &           � � �� o     ����tr  ��      o     �� ���        ���� � �����  �  �         ����
  ' (           � � �� p     �����s  ,�      o     �� ���        ���� � �����  �  �         ����
  ) *           � � �� q     ����Du  t�   ��  o     �� ���       ���� � �����  �  �         ����
  + ,           � � �� r     �����v  �   ��  o     �� ���       ���� � �����  �  �         ����
  - .           � �� s     ����x     ��  o     �� ���       ���� � �����  �  �         ����
  / 0           � 	�� t     ����|y  L+   ��  o     �� ���       ����  �����  �  �         ����
  1 2           � �� u     �����z  �=   ��  o     �� ���       ���� �����  �  �         ����
  3 4           � �� v     ����L|  �O   ��  o     �� ���       ���� �����  �  �         ����
  5 6           � �� w     �����}  $b   ��  o	     �� ���       ���� �����  �  �           ��  # $           � � �� �     ����|o  L�       �       �    �        ���� � �����  �  �           ��  % &           � � �� �     �����p  ��       �      �    �        ���� � �����  �  �           ��  ' (           �  �� �     ����Lr  ��       �      �    �        ���� � �����  �  �         ! ��  ) *           � �� �     �����s  $�       �      �    �        ���� � �����  �  �         ! ��  + ,           � �� �     ����u  l�       �      �    �        ���� � �����  �  �         ! ��  - .           � �� �     �����v  �       �      �    �        ���� � �����  �  �         " ��  / 0           � �� �     �����w  �       �      �    �        ����  �����  �  �         " ��  1 2           � �� �     ����Ty  D)       �      �    �        ���� �����  �  �         " ��  3 4           � $�� �     �����z  �;       �      �    �        ���� �����  �  �         # ��  5 6           � *�� �     ����$|  �M       � 	     �    �        ���� �����  �  �         ����  # $           � � �� n     �����u  ��      }      �� ���        ���� � �����  �  �         ����  % &           �  �� o     ����$w  �      }     �� ���        ���� � �����  �  �         ����  ' (           � �� p     �����x        }     �� ���        ���� � �����  �  �         ����  ) *           � �� q     �����y  d1   ��  }     �� ���       ���� � �����  �  �         ����  + ,           � �� r     ����\{  �C   ��  }     �� ���       ���� � �����  �  �         ����  - .           � �� s     �����|  �U   ��  }     �� ���       ���� � �����  �  �         ����  / 0           � �� t     ����,~  <h   ��  }     �� ���       ����  �����  �  �         ����  1 2           � $�� u     �����  �z   ��  }     �� ���       ���� �����  �  �         ����  3 4           � *�� v     ������  ̌   ��  }     �� ���       ���� �����  �  �         ����  5 6           � 0�� w     ����d�  �   ��  }	     �� ���       ���� �����  �  �         ����	  # $           � � �� n     �����r  ��            �� ���        ���� � �����  �  �         ����	  % &           � � �� o     ����t  4�           �� ���        ���� � �����  �  �         ����	  ' (           � � �� p     ����lu  |�           �� ���        ���� � �����  �  �         ����	  ) *           � � �� q     �����v  �   ��       �� ���       ���� � �����  �  �         ����	  + ,           � � �� r     ����<x     ��       �� ���       ���� � �����  �  �         ����	  - .           � � �� s     �����y  T-   ��       �� ���       ���� � �����  �  �         ����	  / 0           �  �� t     ����{  �?   ��       �� ���       ����  �����  �  �         ����	  1 2           � �� u     ����t|  �Q   ��       �� ���       ���� �����  �  �         ����	  3 4           � �� v     �����}  ,d   ��       �� ���       ���� �����  �  �         ����	  5 6           � �� w     ����D  tv   ��  	     �� ���       ���� �����  �  �         ����  # $           � � �� n     ����,t  <�      #      �� ���        ���� � �����  �  �         ����  % &           � � �� o     �����u  ��      #     �� ���        ���� � �����  �  �         ����  ' (           � �� p     �����v  �
      #     �� ���        ���� � �����  �  �         ����  ) *           � 	�� q     ����dx     ��  #     �� ���       ���� � �����  �  �         ����  + ,           � �� r     �����y  \/   ��  #     �� ���       ���� � �����  �  �         ����  - .           � �� s     ����4{  �A   ��  #     �� ���       ���� � �����  �  �         ����  / 0           � �� t     �����|  �S   ��  #     �� ���       ����  �����  �  �         ����  1 2           � !�� u     ����~  4f   ��  #     �� ���       ���� �����  �  �         ����  3 4           � '�� v     ����l  |x   ��  #     �� ���       ���� �����  �  �         ����  5 6           � -�� w     ����Ԁ  Ċ   ��  #	     �� ���       ���� �����  �  �            ���a�s2    Q�n     �%  $�  ��                 �    ������� � �����  �  �            ���{��2    Z�o     &  "�  d�                �    ������� � �����  �  �            �����2    c�p     \&   �  @�                �    ������� � �����  �  �            ���'�2    l�#q     �&  �                    �   ������� � �����  �  �            ��+�C�2    u�)r     '  �  �C   ��            �   ������� � �����  �  �            ��C�_2    ~�/#s     p'  �  �g   ��            �   ������� � �����  �  �            ��[�{!2    ��5)t     �'  �  ��   ��            �   ������� � �����  �  �            ��s�>2    ��;/u     '(  �  ��   ��            �   ������� � �����  �  �            ���1�[2    ��A5v     �(  �  h�   ��            �   ������� �����  �  �            ���K�x2    ��G;w     �(  �  D�   ��   	         �   �������    �  �  �            ��a�=�2    `�n     �%  �  h�      (       &   �    ������� � �����  �  �            ��T�2    i�o     ,&  �  D�      (      &   �    ������� � �����  �  �            ���5k2    r�p     �&  �         (      &   �    ������� � �����  �  �            ���T�/2    {�#q     �&  �  �0       (      &   �   ������� � �����  �  �            ���s�G2    ��)r     ?'  �  �T   ��  (      &   �   ������� � �����  �  �            �����_2    ��/#s     �'  
�  �x   ��  (      &   �   ������� � �����  �  �            ����w2    ��5)t     �'  �  ��   ��  (      &   �   ������� � �����  �  �            ��3���2    ��;/u     S(  �  l�   ��  (      &   �   ������� � �����  �  �            ��Q���2    ��A5v     �(  �  H�   ��  (      &   �   ������� �����  �  �            ��o�2    ��G;w     
)  �  $   ��  ( 	     &   �   ������� G   �  �  �            ��Y�Y�2    n     �%  `�  ��      <       :   �    ������� � �����  �  �            ��ss2    o     &  ^�  ��      <      :   �    ������� � �����  �  �            ���/�/2    #%#p     g&  \�  x       <      :   �    ������� � �����  �  �            ���J�J2    +++q     �&  Z�  T$       <      :   �   ������� � �����  �  �            ���e�e2    313%r     '  X�  0H   ��  <      :   �   ������� � �����  �  �            ������2    ;7;+s     {'  V�  l   ��  <      :   �   ������� � �����  �  �            ������2    C=C1t     �'  T�  �   ��  <      :   �   ������� � �����  �  �            ����2    KCK7u     2(  R�  ĳ   ��  <      :   �   ������� � �����  �  �            ��)�)�2    SIS=v     �(  P�  ��   ��  <      :   �   ������� �����  �  �            ��C�C�2    [O[Cw     �(  N�  |�   ��  < 	     :   �   ������� y   �  �  �            ���s�a2    [�n     �%  ��  0�      R       O   �    �ؓ���� � �����  �  �            �����{2    d�o     !&  ��  �      R      O   �    �ؓ���� � �����  �  �            �����2    m�p     }&  ��  �      R      O   �    �ؓ���� � �����  �  �            ��'��2    v�#q     �&  ��  �,       R      O   �   �ؓ���� � �����  �  �            ��C�+�2    �)r     4'  ��  �P   ��  R      O   �   �ؓ���� � �����  �  �            ��_C�2    ��/#s     �'  ��  |t   ��  R      O   �   �ؓ���� � �����  �  �            ��{![�2    ��5)t     �'  ��  X�   ��  R      O   �   �ؓ���� � �����  �  �            ���>s2    ��;/u     H(  ��  4�   ��  R      O   �   �ؓ���� � �����  �  �            ���[�12    ��A5v     �(  ��  �   ��  R      O   �   �ؓ���� �����  �  �            ���x�K2    ��G;w     �(  ��  �   ��  R 	     O   �   �ؓ���� �   �  �  �            ��=�a�2    ,�Vn     �%  ��  P�      h       d   �    ��X���� � �����  �  �            ��T�2    2�_o     �%  ��  ,�      h      d   �    ��X���� � �����  �  �            ��k�52    8�hp     R&  ��  �      h      d   �    ��X���� � �����  �  �            ���/�T2    >�qq     �&  ��  �       h      d   �   ��X���� � �����  �  �            ���G�s2    D�z#r     	'  ��  �?   ��  h      d   �   ��X���� � �����  �  �            ���_��2    J��)s     e'  ��  �c   ��  h      d   �   ��X���� � �����  �  �            ���w�2    P��/t     �'  ��  x�   ��  h      d   �   ��X���� � �����  �  �            ����3�2    V��5u     (  ��  T�   ��  h      d   �   ��X���� � �����  �  �            ����Q�2    \��;v     x(  ��  0�   ��  h      d   �   ��X���� �����  �  �            ���o2    b��Aw     �(  ��  �   ��  h 	     d   �   ��X���� �   �  �  �             ��
2    n     �%  ��  ��      �       |   �    ������� � �����  �  �             !�!�
2    o     &  ��  ��      �      |   �    ������� � �����  �  �             :�:�
2    !%#p     r&  ��  �      �      |   �    ������� � �����  �  �             S�S�
2    )++q     �&  ��  �(       �      |   �   ������� � �����  �  �             l
l

2    113%r     *'  ��  hL   ��  �      |   �   ������� � �����  �  �             �%�%
2    97;+s     �'  ��  Dp   ��  �      |   �   ������� � �����  �  �             �@�@
2    A=C1t     �'  ��   �   ��  �      |   �   ������� � �����  �  �             �[�[
2    ICK7u     =(  ��  ��   ��  �      |   �   ������� � �����  �  �             �v�v
2    QIS=v     �(  ��  ��   ��  �      |   �   ������� �����  �  �             ����
2    YO[Cw     �(  ��  ��   ��  � 	     |   �   �������   �  �  �             X��X2    �� � d     �  ��  �T      �       �   �    ������� � �����  �  �             s�o2    �
� � e     �  ��  �t      �      �   �    ������� � �����  �  �             �5��2    �� � f     5   t�  ��      �      �   �    ������� � �����  �  �             �Q�2    �� g     �   T�  ��      �      �   �   ������� � �����  �  �             �m�2    �"
� h     �   4�  t�      �      �   �   ������� � �����  �  �             ��0�2    �*i     )!  �  T�   ��  �      �   �   ������� � �����  �  �             ��E�2    �2
j     {!  ��  4   ��  �      �   �   ������� � �����  �  �             �Z�2    �:k     �!  ��  4   ��  �      �   �   ������� � �����  �  �             0�o2    �B"l     "  ��  �S   ��  �      �   �   ������� �����  �  �             K��'2    �J(m     p"  ��  �s   ��  � 	     �   �   �������    �  �  �             
�=�2    �/n     �%  �  h�      �       �   �    ������� � �����  �  �             '�T�2    �7o     ,&  �  D�      �      �   �    ������� � �����  �  �             D�k2    �?p     �&  �         �      �   �    ������� � �����  �  �             a�/2    �G#q     �&  �  �0       �      �   �   ������� � �����  �  �             ~6�G2    �O)r     ?'  �  �T   ��  �      �   �   ������� � �����  �  �             �T�_2    �W/#s     �'  
�  �x   ��  �      �   �   ������� � �����  �  �             �r�w2    �_5)t     �'  �  ��   ��  �      �   �   ������� � �����  �  �             ����2    �g;/u     S(  �  l�   ��  �      �   �   ������� � �����  �  �             ����2    �oA5v     �(  �  H�   ��  �      �   �   ������� �����  �  �             ��2    wG;w     
)  �  $   ��  � 	     �   �   �������    �  �  �         ����   2 3          d �           	      �        u        ���        ����c   �������������         ����   4 5          g �              >  |        u       ���        ����c   �������������         ����   6 7          j �              \  �        u       ���        ����c   �������������         ����   8 9          m �              z  �        u       ���       ����c   �������������         ����   : ;          p �              �  0        u       ���       ����c   �������������         ����   < =          s �              �  l        u       ���       ����c   �������������         ����   > ?          v �              �  �        u       ���       ����c   �������������         ����   @ A          y �              �  �        u       ���       ����c   �������������         ����   B C          | �                         u       ���       ����c   �������������         ����   D E           �              .  \        u	       ���       ����c   �������������         ����  2 3          d �              �   �         C        ���        ����c   �������������         ����  4 5          g �              �   �        C       ���        ����c   �������������         ����  6 7          j �                        C       ���        ����c   �������������         ����  8 9          m �              "  D        C       ���       ����c   �������������         ����  : ;          p �              @  �        C       ���       ����c   �������������         ����  < =          s �              ^  �        C       ���       ����c   �������������         ����  > ?          v �              |  �        C       ���       ����c   �������������         ����  @ A          y �              �  4        C       ���       ����c   �������������         ����  B C          | �              �  p        C       ���       ����c   �������������         ����  D E           �           	   �  �        C	       ���       ����c   �������������         ����  2 3          d �              ,  h        �        ���        ����c   �������������         ����  4 5          g �              J  �        �       ���        ����c   �������������         ����  6 7          j �              h  �        �       ���        ����c   �������������         ����  8 9          m �              �          �       ���       ����c   �������������         ����  : ;          p �              �  H        �       ���       ����c   �������������         ����  < =          s �           	   �  �        �       ���       ����c   �������������         ����  > ?          v �           	   �  �        �       ���       ����c   �������������         ����  @ A          y �           
   �  �        �       ���       ����c   �������������         ����  B C          | �           
     8        �       ���       ����c   �������������         ����  D E           �              :  t        �	       ���       ����c   �������������         ����  2 3          d �           !   �  /        �        ���        ����c   �������������         ����  4 5          g �           (   �  �        �       ���        ����c   �������������         ����  6 7          j �           )             �       ���        ����c   �������������         ����  8 9          m �           )   *  T        �       ���       ����c   �������������         ����  : ;          p �           *   H  �        �       ���       ����c   �������������         ����  < =          s �           +   f  �        �       ���       ����c   �������������         ����  > ?          v �           +   �          �       ���       ����c   �������������         ����  @ A          y �           ,   �  D        �       ���       ����c   �������������         ����  B C          | �           ,   �  �        �       ���       ����c   �������������         ����  D E           �           -   �  �        �	       ���       ����c   �������������         ����  3 4          d �              �  F        u        ���        ����c   �������������         ����  5 6          g �              �  �	        u       ���        ����c   �������������         ����  7 8          j �              �  �	        u       ���        ����c   �������������         ����  9 :          m �              
  
        u       ���       ����c   �������������         ����  ; <          p �              (  P
        u       ���       ����c   �������������         ����  = >          s �              F  �
        u       ���       ����c   �������������         ����  ? @          v �              d  �
        u       ���       ����c   �������������         ����  A B          y �              �          u       ���       ����c   �������������         ����  C D          | �              �  @        u       ���       ����c   �������������         ����  E F           �              �  |        u	       ���       ����c   �������������         ����  4 5          d �              @  �                ���        ����c   �������������         ����  6 7          g �               ^  �               ���        ����c   �������������         ����  8 9          j �           !   |  �               ���        ����c   �������������         ����  : ;          m �           !   �  4               ���       ����c   �������������         ����  < =          p �           "   �  p               ���       ����c   �������������         ����  > ?          s �           #   �  �               ���       ����c   �������������         ����  @ A          v �           #   �  �               ���       ����c   �������������         ����  B C          y �           $     $               ���       ����c   �������������         ����  D E          | �           $   0  `               ���       ����c   �������������         ����  F G           �           %   N  �        	       ���       ����c   �������������             �@U�2    K K              �  �        �       �   �    �������c   �������������             �BW�2    P K                        �      �   �    �������c   �������������             �DY�2    U K                 @        �      �   �    �������c   �������������             �F[�2    Z K              >  |        �      �   �   �������c   �������������             �H]�2    _ K              \  �        �      �   �   �������c   �������������             �J_�2    d K              z  �        �      �   �   �������c   �������������             �La�2    i K              �  0        �      �   �   �������c   �������������             �Nc�2    n K              �  l        �      �   �   �������c   �������������             �Pe�2    s K              �  �        �      �   �   �������c   �������������             �Rg�2    x K              �  �        � 	     �   �   �������c   �������������          ��  r  D F x d     U d           �   �  �        �       ��	 ���        ������  ����������������        ��  r  � � x d (    �           �   X          �       ��	 ���        ������  ����������������       ��  r  PRx d <    GS         �      �        �       ��	 ���        ������  ����������������       ��  r  ��x d P    ��E        �   L  |        �       ��	 ���        ������  ����������������       ��  r  \^x d d    ��O O       �   �  (#        �       ��	 ��         ������  ����������������        ��t ��                           ������  �      M      �� ��        ������  ����������������        ��t ��                           ���� � @B      N      �� ��        ������  ����������������        ��t ��                           ����@B ��      O      �� ��        ������  ����������������        ��t ��                           ������  �      P      �� ��        ������  ����������������        ��t ��                           ���� � @B      Q      �� ��        ������  ����������������        ��t ��                           ����@B ��      R      �� ��        ������  ����������������        ��t ��                           ������  �      S      �� ��        ������  ����������������        ��t ��                           ���� � @B      T      �� ��        ������  ����������������        ��t ��            	               ����@B ��      U      �� ��	        ������  ����������������        ��t ��            
               ���� � @B      V      �� ��
        ������  ����������������        ��t ��                           �����q `�      W      �� ��        ������  ����������������        ��t ��                           ����@B ��      X      �� ��        ������  ����������������       ����� ��                            �����  �       A      ��b ��        ������  ����������������        ��t ��                           ����'   N       Y      �� ��        ������  ����������������       ����u �� 
 ��                    @B  � ��      d      �� ��        ������  ����������������       ����u ��<  ��	                    �� @B  	=      e      �� ��        ������  ����������������       ����u ��Z  ��                    ��- `� ��[      f      �� ��        ������  ����������������       ����u ��
  ��                    @B  � ��      g      �� ��        ������  ����������������       ����u �� < ��	                    �� @B  	=      h      �� ��        ������  ����������������       ����u �� Z ��                    ��- `� ��[      i      �� ��        ������  ����������������       ��  v ��    ��                    @B  � ��      j      �� ��        ������  ����������������       �� v ��    ��	                    �� @B  	=      k      �� ��        ������  ����������������       �� v ��    ��                    ��- `� ��[      l      �� ��        ������  ����������������        ��w ��F F ��	                    @B  � ��      m      �� ��        ������  ����������������          ��Z	�92    ��0$x     �,  
�  �q                     ������� � �����  �  �            ��t$�X2    ��6*y     -  &�  ҙ                    ������� � �����  �  �            ���?�w2    ��<0z     u-  B�  ��   ��                ������� � �����  �  �            ���Z��2    ��B6{     �-  ^�  ��   ��               ������� � �����  �  �            ���u��2    ��H<|     B.  z�     ��               ������� � �����  �  �            �����2    ��NB}     �.  ��  ":   ��               ������� � �����  �  �            ����8�2    ��TH~     /  ��  6b   ��               ������� � �����  �  �            ���U2    ��ZN     v/  ��  J�   ��               ������� �����  �  �            ��*�r12    �`T�     �/  ��  ^�   ��               ������� �����  �  �            ��D��P2    �fZ�     C0  �  r�   ��   	            ������� 
   �  �  �            ��,��{2    ��0$x     �,  ��  ��      )       '       ������� � �����  �  �            ��K���2    ��6*y     <-  �  ��      )      '       ������� � �����  �  �            ��j��2    ��<0z     �-  2�  ��   ��  )      '       ������� � �����  �  �            ���4
�2    ��B6{     	.  N�  ��   ��  )      '      ������� � �����  �  �            ���U"�2    ��H<|     p.  j�  �#   ��  )      '      ������� � �����  �  �            ���v:�2    ��NB}     �.  ��  �K   ��  )      '      ������� � �����  �  �            ����R2    �TH~     =/  ��  t   ��  )      '      ������� � �����  �  �            ���j*2    �ZN     �/  ��  �   ��  )      '      ������� �����  �  �            ��$��C2    �`T�     
0  ��  .�   ��  )      '      ������� �����  �  �            ��C��\2    �fZ�     q0  ��  B�   ��  ) 	     '      ������� 
Q   �  �  �            ������2    ?8?,x     �,  F�  2v      =       ;       ������� � �����  �  �            ����2    G>G2y     -  b�  F�      =      ;       ������� � �����  �  �            ��4�4�2    ODO8z     �-  ~�  Z�   ��  =      ;       ������� � �����  �  �            ��PP2    WJW>{     �-  ��  n�   ��  =      ;      ������� � �����  �  �            ��ll2    _P_D|     N.  ��  �   ��  =      ;      ������� � �����  �  �            ���<�<2    gVgJ}     �.  ��  �>   ��  =      ;      ������� � �����  �  �            ���Y�Y2    o\oP~     /  ��  �f   ��  =      ;      ������� � �����  �  �            ���v�v2    wbwV     �/  
�  ��   ��  =      ;      ������� �����  �  �            ������2    h\�     �/  &�  Ҷ   ��  =      ;      ������� �����  �  �            ������2    �n�b�     O0  B�  ��   ��  = 	     ;      ������� 
�   �  �  �            ���9Z	2    ��0$x     �,  ��        S       P       ������� � �����  �  �            ���Xt$2    ��6*y     1-  ��  .�      S      P       ������� � �����  �  �            ���w�?2    ��<0z     �-  ��  B�   ��  S      P       ������� � �����  �  �            �����Z2    ��B6{     �-  �  V�   ��  S      P      ������� � �����  �  �            �����u2    ��H<|     d.  .�  j   ��  S      P      ������� � �����  �  �            �����2    ��NB}     �.  J�  ~G   ��  S      P      ������� � �����  �  �            ��8���2    �TH~     2/  f�  �o   ��  S      P      ������� � �����  �  �            ��U�2    �	ZN     �/  ��  ��   ��  S      P      ������� �����  �  �            ��r1*�2    �`T�     �/  ��  ��   ��  S      P      ������� �����  �  �            ���PD�2    �fZ�     e0  ��  ��   ��  S 	     P      ������� 
�   �  �  �            ���{,�2    K��*x     �,  ��  Jm      i       e       ������� � �����  �  �            ����K�2    R��0y     -  ��  ^�      i      e       ������� � �����  �  �            ����j2    Y��6z     j-  �  r�   ��  i      e       ������� � �����  �  �            ��
��42    `��<{     �-  "�  ��   ��  i      e      ������� � �����  �  �            ��"��U2    g��B|     7.  >�  �   ��  i      e      ������� � �����  �  �            ��:��v2    n��H}     �.  Z�  �5   ��  i      e      ������� � �����  �  �            ��R��2    u��N~     /  v�  �]   ��  i      e      ������� � �����  �  �            ��j*�2    |��T     k/  ��  օ   ��  i      e      ������� �����  �  �            ���C$�2    ���Z�     �/  ��  �   ��  i      e      ������� �����  �  �            ���\C�2    ���`�     80  ��  ��   ��  i 	     e      ������� 
�   �  �  �             �P�P
2    =8?,x     �,  ��  �z      �       }       ������� � �����  �  �             �l�l
2    E>G2y     %-  ��  ��      �      }       ������� � �����  �  �             ����
2    MDO8z     �-  ��  ��   ��  �      }       ������� � �����  �  �             ����
2    UJW>{     �-  ��  ��   ��  �      }      ������� � �����  �  �             ��
2    ]P_D|     Y.  ��  �   ��  �      }      ������� � �����  �  �             (�(�
2    eVgJ}     �.  �  
C   ��  �      }      ������� � �����  �  �             C�C�
2    m\oP~     &/  *�  k   ��  �      }      ������� � �����  �  �             ^^
2    ubwV     �/  F�  2�   ��  �      }      ������� �����  �  �             y0y0
2    }h\�     �/  b�  F�   ��  �      }      ������� �����  �  �             �L�L
2    �n�b�     Z0  ~�  Z�   ��  � 	     }      ������� 
  �  �  �             ���{2    �[0$x     �,  ��  ��      �       �       ������� � �����  �  �             ����2    �d6*y     <-  �  ��      �      �       ������� � �����  �  �             ���2    �m<0z     �-  2�  ��   ��  �      �       ������� � �����  �  �             %�
�2    �vB6{     	.  N�  ��   ��  �      �      ������� � �����  �  �             C"�2    H<|     p.  j�  �#   ��  �      �      ������� � �����  �  �             a.:�2    �NB}     �.  ��  �K   ��  �      �      ������� � �����  �  �             NR2    �TH~     =/  ��  t   ��  �      �      ������� � �����  �  �             �nj*2    �ZN     �/  ��  �   ��  �      �      ������� �����  �  �             ���C2    %�`T�     
0  ��  .�   ��  �      �      ������� �����  �  �             ���\2    -�fZ�     q0  ��  B�   ��  � 	     �      ������� 
   �  �  �         ����x ��                                        /     n      ��L ��        ������  ����������������       ����x ��                                       /     o      ��M ��        ������  ����������������       ����x ��                                       /     p      ��N ��        ������  ����������������       ����x ��                                       /     q      ��O ��        ������  ����������������       ����� ��                            �����  �        B      ��c ��        ������  ����������������        ��j ��          ^               ����'  �#        
      ��c ��        ������  ����������������        ��p ��  3                        �����  �        8      ��c ��        ������  ����������������        ��p ��  9                        �����  �        9      ��c ��         ������  ����������������        ��p ��  ?                        �����  �        :      ��c ��!        ������  ����������������        ��p ��  ,                        �����  �        ;      ��c ��"        ������  ����������������        ��p ��  N                        �����  �        <      ��c ��#        ������  ����������������        ��p ��  j                        �����  �        =      ��c ��$        ������  ����������������       ����� ��                            �����  �        C      ��d ��%        ������  ����������������       ����� ��                            �����  �        D      ��d ��%        ������  ����������������       ����� ��                            �����  �        E      ��d ��%        ������  ����������������       ����� ��                            �����  �        F      ��d ��%        ������  ����������������        ��t ��                           ����'   N       Z      �� ��&        ������  ����������������        ��t ��                           ����'   N       [      �� ��&        ������  ����������������        ��t ��                           ����'   N       \      �� ��&        ������  ����������������        ��t ��                           ����'   N       ]      �� ��&        ������  ����������������       ����   A B          �� � x       �y  X�      "        ��'        ���� � �����  �  �         ����   C D          �� � y     I  z{  ��       "       ��'        ���� � �����  �  �         ����   E F          �$� � z     �   }   �   ��  "       ��'        ���� � �����  �  �         ����   H I          �*� � {     �  �~  T�   ��  "       ��'       ���� � �����  �  �         ����   J K          �0� � |     �  �  �    ��  "       ��'       ����  �����  �  �         ����   L M          �6� � }     #  ��  �   ��  "       ��'       ���� �����  �  �         ����   N O          <� � ~     Z  �  P+   ��  "       ��'       ���� �����  �  �         ����   P Q          B� �      �  ��  �@   ��  "       ��'       ���� �����  �  �         ����   S T          H� � �     �  $�  �U   ��  "       ��'       ���� �����  �  �         ����   U V          N� � �     �  ��  Lk   ��  "	       ��'       ���� #K  �  �  �         ����   3 4          � �� x       �y  X�      6        ��(        ���� � �����  �  �         ����   5 6          � �� y     I  z{  ��       6       ��(        ���� � �����  �  �         ����   7 8          � !�� z     �   }   �   ��  6       ��(        ���� � �����  �  �         ����   9 :          � '�� {     �  �~  T�   ��  6       ��(       ���� � �����  �  �         ����   ; <          � -�� |     �  �  �    ��  6       ��(       ����  �����  �  �         ����   = >          � 3�� }     #  ��  �   ��  6       ��(       ���� �����  �  �         ����   @ A          � 9�� ~     Z  �  P+   ��  6       ��(       ���� �����  �  �         ����   B C          � ?�      �  ��  �@   ��  6       ��(       ���� �����  �  �         ����   D E          � E� �     �  $�  �U   ��  6       ��(       ���� �����  �  �         ����   F G          � K� �     �  ��  Lk   ��  6	       ��(       ���� #K  �  �  �         ����   2 3          �� �� x       �y  X�      J        ��)        ���� � �����  �  �         ����   4 5          �� �� y     I  z{  ��       J       ��)        ���� � �����  �  �         ����   6 7          �� �� z     �   }   �   ��  J       ��)        ���� � �����  �  �         ����   8 9          �� �� {     �  �~  T�   ��  J       ��)       ���� � �����  �  �         ����   : ;          �� �� |     �  �  �    ��  J       ��)       ����  �����  �  �         ����   < =          �� �� }     #  ��  �   ��  J       ��)       ���� �����  �  �         ����   ? @          �� �� ~     Z  �  P+   ��  J       ��)       ���� �����  �  �         ����   A B          �� ��      �  ��  �@   ��  J       ��)       ���� �����  �  �         ����   C D          �� �� �     �  $�  �U   ��  J       ��)       ���� �����  �  �         ����   E F          �� �� �     �  ��  Lk   ��  J	       ��)       ���� #K  �  �  �         ����   & '          � 
�� x       �y  X�      ^        ��*        ���� � �����  �  �         ����   ( )          � �� y     I  z{  ��       ^       ��*        ���� � �����  �  �         ����   * +          � �� z     �   }   �   ��  ^       ��*        ���� � �����  �  �         ����   , -          � �� {     �  �~  T�   ��  ^       ��*       ���� � �����  �  �         ����   . /          � "�� |     �  �  �    ��  ^       ��*       ����  �����  �  �         ����   0 1          � (�� }     #  ��  �   ��  ^       ��*       ���� �����  �  �         ����   2 3          � .� ~     Z  �  P+   ��  ^       ��*       ���� �����  �  �         ����   4 5          � 4	�      �  ��  �@   ��  ^       ��*       ���� �����  �  �         ����   6 7          � :� �     �  $�  �U   ��  ^       ��*       ���� �����  �  �         ����   8 9          � @� �     �  ��  Lk   ��  ^	       ��*       ���� #K  �  �  �         ����   3 4          hn� � x       �y  X�      r        ��+        ���� � �����  �  �         ����   5 6          ou� � y     I  z{  ��       r       ��+        ���� � �����  �  �         ����   7 8          v|� � z     �   }   �   ��  r       ��+        ���� � �����  �  �         ����   9 :          }�� � {     �  �~  T�   ��  r       ��+       ���� � �����  �  �         ����   ; <          ��� � |     �  �  �    ��  r       ��+       ����  �����  �  �         ����   = >          ��� � }     #  ��  �   ��  r       ��+       ���� �����  �  �         ����   @ A          ��� � ~     Z  �  P+   ��  r       ��+       ���� �����  �  �         ����   B C          ��� �      �  ��  �@   ��  r       ��+       ���� �����  �  �         ����   D E          ��� � �     �  $�  �U   ��  r       ��+       ���� �����  �  �         ����   F G          ��� � �     �  ��  Lk   ��  r	       ��+       ���� #K  �  �  �         ����  ? @          �� � x     �   x   �      �        ��,        ���� � �����  �  �         ����  A B          �� � y       �y  T�       �       ��,        ���� � �����  �  �         ����  C D          �$� � z     :  {  ��   ��  �       ��,        ���� � �����  �  �         ����  F G          �*� � {     p  �|  ��   ��  �       ��,       ���� � �����  �  �         ����  H I          �0� � |     �  ~  P�   ��  �       ��,       ����  �����  �  �         ����  J K          �6� � }     �  �  ��   ��  �       ��,       ���� �����  �  �         ����  L M          �<� � ~       $�  �   ��  �       ��,       ���� �����  �  �         ����  N O          �B� �      K  ��  L%   ��  �       ��,       ���� �����  �  �         ����  Q R          H� � �     �  0�  �:   ��  �       ��,       ���� �����  �  �         ����  S T          	N� � �     �  ��  �O   ��  �	       ��,       ���� #K  �  �  �         ����  2 3          �  �� x     �   x   �      �        ��-        ���� � �����  �  �         ����  4 5          � �� y       �y  T�       �       ��-        ���� � �����  �  �         ����  6 7          � �� z     :  {  ��   ��  �       ��-        ���� � �����  �  �         ����  8 9          � �� {     p  �|  ��   ��  �       ��-       ���� � �����  �  �         ����  : ;          � �� |     �  ~  P�   ��  �       ��-       ����  �����  �  �         ����  < =          � �� }     �  �  ��   ��  �       ��-       ���� �����  �  �         ����  ? @          � $�� ~       $�  �   ��  �       ��-       ���� �����  �  �         ����  A B          � *��      K  ��  L%   ��  �       ��-       ���� �����  �  �         ����  C D          � 0�� �     �  0�  �:   ��  �       ��-       ���� �����  �  �         ����  E F          � 6� �     �  ��  �O   ��  �	       ��-       ���� #K  �  �  �         ����  1 2          o� o� x     �   x   �      �        ��.        ���� � �����  �  �         ����  3 4          v� v� y       �y  T�       �       ��.        ���� � �����  �  �         ����  5 6          }� }� z     :  {  ��   ��  �       ��.        ���� � �����  �  �         ����  7 8          �� �� {     p  �|  ��   ��  �       ��.       ���� � �����  �  �         ����  9 :          �� �� |     �  ~  P�   ��  �       ��.       ����  �����  �  �         ����  ; <          �� �� }     �  �  ��   ��  �       ��.       ���� �����  �  �         ����  > ?          �� �� ~       $�  �   ��  �       ��.       ���� �����  �  �         ����  @ A          �� ��      K  ��  L%   ��  �       ��.       ���� �����  �  �         ����  B C          �� �� �     �  0�  �:   ��  �       ��.       ���� �����  �  �         ����  D E          �� �� �     �  ��  �O   ��  �	       ��.       ���� #K  �  �  �         ����  % &          � �� x     �   x   �      �        ��/        ���� � �����  �  �         ����  ' (          � �� y       �y  T�       �       ��/        ���� � �����  �  �         ����  ) *          � �� z     :  {  ��   ��  �       ��/        ���� � �����  �  �         ����  + ,          � �� {     p  �|  ��   ��  �       ��/       ���� � �����  �  �         ����  - .          � �� |     �  ~  P�   ��  �       ��/       ����  �����  �  �         ����  / 0          � �� }     �  �  ��   ��  �       ��/       ���� �����  �  �         ����  1 2          � %�� ~       $�  �   ��  �       ��/       ���� �����  �  �         ����  3 4          � + �      K  ��  L%   ��  �       ��/       ���� �����  �  �         ����  5 6          � 1� �     �  0�  �:   ��  �       ��/       ���� �����  �  �         ����  7 8          � 7� �     �  ��  �O   ��  �	       ��/       ���� #K  �  �  �         ����  3 4          hd� � x     �   x   �      �        ��0        ���� � �����  �  �         ����  5 6          ok� � y       �y  T�       �       ��0        ���� � �����  �  �         ����  7 8          vr� � z     :  {  ��   ��  �       ��0        ���� � �����  �  �         ����  9 :          }y� � {     p  �|  ��   ��  �       ��0       ���� � �����  �  �         ����  ; <          ��� � |     �  ~  P�   ��  �       ��0       ����  �����  �  �         ����  = >          ��� � }     �  �  ��   ��  �       ��0       ���� �����  �  �         ����  @ A          ��� � ~       $�  �   ��  �       ��0       ���� �����  �  �         ����  B C          ��� �      K  ��  L%   ��  �       ��0       ���� �����  �  �         ����  D E          ��� � �     �  0�  �:   ��  �       ��0       ���� �����  �  �         ����  F G          ��� � �     �  ��  �O   ��  �	       ��0       ���� #K  �  �  �         $ ��  B C           �� � �     ����ā  �       �       �    1        ���� � �����  �  �         $ ��  D E           �� � �     ����J�  .       �      �    1        ���� � �����  �  �         $ ��  F G           �$� � �     ����Є  `C       �      �    1        ���� � �����  �  �         $ ��  I J            *� � �     ����V�  �X       �      �    1        ���� � �����  �  �         $ ��  K L           0� � �     ����܇  n       �      �    1        ����  �����  �  �         $ ��  M N           6� � �     ����b�  \�       �      �    1        ���� �����  �  �         $ ��  O P           <� � �     �����  ��       �      �    1        ���� �����  �  �         $ ��  Q R            B� � �     ����n�  �       �      �    1        ���� �����  �  �         $ ��  T U           (H� � �     �����  X�       �      �    1        ���� �����  �  �         $ ��  V W           0N� � �     ����z�  ��       � 	     �    1        ���� #�����  �  �         $ ��  3 4           � '�� �     ����ā  �       �       �    1        ���� � �����  �  �         $ ��  5 6           � -�� �     ����J�  .       �      �    1        ���� � �����  �  �         $ ��  7 8           � 3�� �     ����Є  `C       �      �    1        ���� � �����  �  �         $ ��  9 :           � 9�� �     ����V�  �X       �      �    1        ���� � �����  �  �         $ ��  ; <           � ?� �     ����܇  n       �      �    1        ����  �����  �  �         $ ��  = >           � E	� �     ����b�  \�       �      �    1        ���� �����  �  �         $ ��  @ A           � K� �     �����  ��       �      �    1        ���� �����  �  �         $ ��  B C           Q� �     ����n�  �       �      �    1        ���� �����  �  �         $ ��  D E           W!� �     �����  X�       �      �    1        ���� �����  �  �         $ ��  F G           ])� �     ����z�  ��       � 	     �    1        ���� #�����  �  �         $ ��  2 3           �� �� �     ����ā  �       �       �    1        ���� � �����  �  �         $ ��  4 5           �� �� �     ����J�  .       �      �    1        ���� � �����  �  �         $ ��  6 7           �� �� �     ����Є  `C       �      �    1        ���� � �����  �  �         $ ��  8 9           �� �� �     ����V�  �X       �      �    1        ���� � �����  �  �         $ ��  : ;           �� �� �     ����܇  n       �      �    1        ����  �����  �  �         $ ��  < =           �� �� �     ����b�  \�       �      �    1        ���� �����  �  �         $ ��  ? @           �� �� �     �����  ��       �      �    1        ���� �����  �  �         $ ��  A B           �� �� �     ����n�  �       �      �    1        ���� �����  �  �         $ ��  C D           �� �� �     �����  X�       �      �    1        ���� �����  �  �         $ ��  E F           �� �� �     ����z�  ��       � 	     �    1        ���� #�����  �  �         $ ��  & '           � �� �     ����ā  �       �       �    1        ���� � �����  �  �         $ ��  ( )           � �� �     ����J�  .       �      �    1        ���� � �����  �  �         $ ��  * +           � �� �     ����Є  `C       �      �    1        ���� � �����  �  �         $ ��  , -           � $�� �     ����V�  �X       �      �    1        ���� � �����  �  �         $ ��  . /           � *�� �     ����܇  n       �      �    1        ����  �����  �  �         $ ��  0 1           � 0�� �     ����b�  \�       �      �    1        ���� �����  �  �         $ ��  2 3           � 6� �     �����  ��       �      �    1        ���� �����  �  �         $ ��  4 5           � <� �     ����n�  �       �      �    1        ���� �����  �  �         $ ��  6 7           � B� �     �����  X�       �      �    1        ���� �����  �  �         $ ��  8 9           � H� �     ����z�  ��       � 	     �    1        ���� #�����  �  �         $ ��  4 5           hy� � �     ����ā  �             �     1        ���� � �����  �  �         $ ��  6 7           o�� � �     ����J�  .            �     1        ���� � �����  �  �         $ ��  8 9           v�� � �     ����Є  `C            �     1        ���� � �����  �  �         $ ��  : ;           }�� � �     ����V�  �X            �     1        ���� � �����  �  �         $ ��  < =           ��� � �     ����܇  n            �     1        ����  �����  �  �         $ ��  > ?           ��� � �     ����b�  \�            �     1        ���� �����  �  �         $ ��  A B           ��� � �     �����  ��            �     1        ���� �����  �  �         $ ��  C D           ��� � �     ����n�  �            �     1        ���� �����  �  �         $ ��  E F           ��� � �     �����  X�            �     1        ���� �����  �  �         $ ��  G H           ��� � �     ����z�  ��       	     �     1        ���� #�����  �  �         ����  @ A          �� � x     �  �w  ��      �        ��2        ���� � �����  �  �         ����  B C          �� � y     �  "y  ܟ       �       ��2        ���� � �����  �  �         ����  D E          �$� � z     ,  �z  0�   ��  �       ��2        ���� � �����  �  �         ����  G H          �*� � {     b  .|  ��   ��  �       ��2       ���� � �����  �  �         ����  I J          �0� � |     �  �}  ��   ��  �       ��2       ����  �����  �  �         ����  K L          �6� � }     �  :  ,�   ��  �       ��2       ���� �����  �  �         ����  M N          �<� � ~       ��  �
   ��  �       ��2       ���� �����  �  �         ����  O P          B� �      =  F�  �   ��  �       ��2       ���� �����  �  �         ����  R S          H� � �     s  ̃  (5   ��  �       ��2       ���� �����  �  �         ����  T U          N� � �     �  R�  |J   ��  �	       ��2       ���� #K  �  �  �         ����  2 3          � �� x     �  �w  ��              ��3        ���� � �����  �  �         ����  4 5          � �� y     �  "y  ܟ              ��3        ���� � �����  �  �         ����  6 7          � �� z     ,  �z  0�   ��         ��3        ���� � �����  �  �         ����  8 9          � �� {     b  .|  ��   ��         ��3       ���� � �����  �  �         ����  : ;          � %�� |     �  �}  ��   ��         ��3       ����  �����  �  �         ����  < =          � +�� }     �  :  ,�   ��         ��3       ���� �����  �  �         ����  ? @          � 1�� ~       ��  �
   ��         ��3       ���� �����  �  �         ����  A B          � 7��      =  F�  �   ��         ��3       ���� �����  �  �         ����  C D          � =� �     s  ̃  (5   ��         ��3       ���� �����  �  �         ����  E F          � C� �     �  R�  |J   ��  	       ��3       ���� #K  �  �  �         ����  1 2          |� |� x     �  �w  ��              ��4        ���� � �����  �  �         ����  3 4          �� �� y     �  "y  ܟ              ��4        ���� � �����  �  �         ����  5 6          �� �� z     ,  �z  0�   ��         ��4        ���� � �����  �  �         ����  7 8          �� �� {     b  .|  ��   ��         ��4       ���� � �����  �  �         ����  9 :          �� �� |     �  �}  ��   ��         ��4       ����  �����  �  �         ����  ; <          �� �� }     �  :  ,�   ��         ��4       ���� �����  �  �         ����  > ?          �� �� ~       ��  �
   ��         ��4       ���� �����  �  �         ����  @ A          �� ��      =  F�  �   ��         ��4       ���� �����  �  �         ����  B C          �� �� �     s  ̃  (5   ��         ��4       ���� �����  �  �         ����  D E          �� �� �     �  R�  |J   ��  	       ��4       ���� #K  �  �  �         ����  % &          � �� x     �  �w  ��      /        ��5        ���� � �����  �  �         ����  ' (          � �� y     �  "y  ܟ       /       ��5        ���� � �����  �  �         ����  ) *          � �� z     ,  �z  0�   ��  /       ��5        ���� � �����  �  �         ����  + ,          � �� {     b  .|  ��   ��  /       ��5       ���� � �����  �  �         ����  - .          � $�� |     �  �}  ��   ��  /       ��5       ����  �����  �  �         ����  / 0          � *�� }     �  :  ,�   ��  /       ��5       ���� �����  �  �         ����  1 2          � 0�� ~       ��  �
   ��  /       ��5       ���� �����  �  �         ����  3 4          � 6�      =  F�  �   ��  /       ��5       ���� �����  �  �         ����  5 6          � <� �     s  ̃  (5   ��  /       ��5       ���� �����  �  �         ����  7 8          � B� �     �  R�  |J   ��  /	       ��5       ���� #K  �  �  �         ����  3 4          hm� � x     �  �w  ��      @        ��6        ���� � �����  �  �         ����  5 6          ot� � y     �  "y  ܟ       @       ��6        ���� � �����  �  �         ����  7 8          v{� � z     ,  �z  0�   ��  @       ��6        ���� � �����  �  �         ����  9 :          }�� � {     b  .|  ��   ��  @       ��6       ���� � �����  �  �         ����  ; <          ��� � |     �  �}  ��   ��  @       ��6       ����  �����  �  �         ����  = >          ��� � }     �  :  ,�   ��  @       ��6       ���� �����  �  �         ����  @ A          ��� � ~       ��  �
   ��  @       ��6       ���� �����  �  �         ����  B C          ��� �      =  F�  �   ��  @       ��6       ���� �����  �  �         ����  D E          ��� � �     s  ̃  (5   ��  @       ��6       ���� �����  �  �         ����  F G          ��� � �     �  R�  |J   ��  @	       ��6       ���� #K  �  �  �         ����  ? @          �� � x     �  �~  ��      b        ��7        ���� � �����  �  �         ����  A B          �� � y     �  *�  L       b       ��7        ���� � �����  �  �         ����  C D          �$� � z     (  ��  �   ��  b       ��7        ���� � �����  �  �         ����  F G          �*� � {     ^  6�  �,   ��  b       ��7       ���� � �����  �  �         ����  H I          �0� � |     �  ��  HB   ��  b       ��7       ����  �����  �  �         ����  J K          �6� � }     �  B�  �W   ��  b       ��7       ���� �����  �  �         ����  L M          �<� � ~       ȇ  �l   ��  b       ��7       ���� �����  �  �         ����  N O          �B� �      9  N�  D�   ��  b       ��7       ���� �����  �  �         ����  Q R          �H� � �     o  Ԋ  ��   ��  b       ��7       ���� �����  �  �         ����  S T          N� � �     �  Z�  �   ��  b	       ��7       ���� #K  �  �  �         ����  2 3          � � �� x     �  �~  ��      s        ��8        ���� � �����  �  �         ����  4 5          � �� y     �  *�  L       s       ��8        ���� � �����  �  �         ����  6 7          � �� z     (  ��  �   ��  s       ��8        ���� � �����  �  �         ����  8 9          � �� {     ^  6�  �,   ��  s       ��8       ���� � �����  �  �         ����  : ;          � �� |     �  ��  HB   ��  s       ��8       ����  �����  �  �         ����  < =          � �� }     �  B�  �W   ��  s       ��8       ���� �����  �  �         ����  ? @          � �� ~       ȇ  �l   ��  s       ��8       ���� �����  �  �         ����  A B          � %��      9  N�  D�   ��  s       ��8       ���� �����  �  �         ����  C D          � +�� �     o  Ԋ  ��   ��  s       ��8       ���� �����  �  �         ����  E F          � 1�� �     �  Z�  �   ��  s	       ��8       ���� #K  �  �  �         ����  1 2          j� j� x     �  �~  ��      �        ��9        ���� � �����  �  �         ����  3 4          q� q� y     �  *�  L       �       ��9        ���� � �����  �  �         ����  5 6          x� x� z     (  ��  �   ��  �       ��9        ���� � �����  �  �         ����  7 8          � � {     ^  6�  �,   ��  �       ��9       ���� � �����  �  �         ����  9 :          �� �� |     �  ��  HB   ��  �       ��9       ����  �����  �  �         ����  ; <          �� �� }     �  B�  �W   ��  �       ��9       ���� �����  �  �         ����  > ?          �� �� ~       ȇ  �l   ��  �       ��9       ���� �����  �  �         ����  @ A          �� ��      9  N�  D�   ��  �       ��9       ���� �����  �  �         ����  B C          �� �� �     o  Ԋ  ��   ��  �       ��9       ���� �����  �  �         ����  D E          �� �� �     �  Z�  �   ��  �	       ��9       ���� #K  �  �  �         ����  % &          � � �� x     �  �~  ��      �        ��:        ���� � �����  �  �         ����  ' (          � �� y     �  *�  L       �       ��:        ���� � �����  �  �         ����  ) *          � 
�� z     (  ��  �   ��  �       ��:        ���� � �����  �  �         ����  + ,          � �� {     ^  6�  �,   ��  �       ��:       ���� � �����  �  �         ����  - .          � �� |     �  ��  HB   ��  �       ��:       ����  �����  �  �         ����  / 0          � �� }     �  B�  �W   ��  �       ��:       ���� �����  �  �         ����  1 2          � "�� ~       ȇ  �l   ��  �       ��:       ���� �����  �  �         ����  3 4          � (��      9  N�  D�   ��  �       ��:       ���� �����  �  �         ����  5 6          � .� �     o  Ԋ  ��   ��  �       ��:       ���� �����  �  �         ����  7 8          � 4� �     �  Z�  �   ��  �	       ��:       ���� #K  �  �  �         ����  3 4          ha� � x     �  �~  ��      �        ��;        ���� � �����  �  �         ����  5 6          oh� � y     �  *�  L       �       ��;        ���� � �����  �  �         ����  7 8          vo� � z     (  ��  �   ��  �       ��;        ���� � �����  �  �         ����  9 :          }v� � {     ^  6�  �,   ��  �       ��;       ���� � �����  �  �         ����  ; <          �}� � |     �  ��  HB   ��  �       ��;       ����  �����  �  �         ����  = >          ��� � }     �  B�  �W   ��  �       ��;       ���� �����  �  �         ����  @ A          ��� � ~       ȇ  �l   ��  �       ��;       ���� �����  �  �         ����  B C          ��� �      9  N�  D�   ��  �       ��;       ���� �����  �  �         ����  D E          ��� � �     o  Ԋ  ��   ��  �       ��;       ���� �����  �  �         ����  F G          ��� � �     �  Z�  �   ��  �	       ��;       ���� #K  �  �  �         ����  B C          �� � x     �  }  �      �        ��<        ���� � �����  �  �         ����  D E          �� � y     �  �~  l�       �       ��<        ���� � �����  �  �         ����  F G          �$� � z     �   �  �   ��  �       ��<        ���� � �����  �  �         ����  I J          �*� � {     &  ��     ��  �       ��<       ���� � �����  �  �         ����  K L          0� � |     ]  ,�  h,   ��  �       ��<       ����  �����  �  �         ����  M N          6� � }     �  ��  �A   ��  �       ��<       ���� �����  �  �         ����  O P          <� � ~     �  8�  W   ��  �       ��<       ���� �����  �  �         ����  Q R          B� �        ��  dl   ��  �       ��<       ���� �����  �  �         ����  T U          #H� � �     7  D�  ��   ��  �       ��<       ���� �����  �  �         ����  V W          +N� � �     n  ʊ  �   ��  �	       ��<       ���� #K  �  �  �         ����  3 4          � "�� x     �  }  �      �        ��=        ���� � �����  �  �         ����  5 6          � (�� y     �  �~  l�       �       ��=        ���� � �����  �  �         ����  7 8          � .�� z     �   �  �   ��  �       ��=        ���� � �����  �  �         ����  9 :          � 4�� {     &  ��     ��  �       ��=       ���� � �����  �  �         ����  ; <          � :�� |     ]  ,�  h,   ��  �       ��=       ����  �����  �  �         ����  = >          � @� }     �  ��  �A   ��  �       ��=       ���� �����  �  �         ����  @ A          � F� ~     �  8�  W   ��  �       ��=       ���� �����  �  �         ����  B C          � L�        ��  dl   ��  �       ��=       ���� �����  �  �         ����  D E          R� �     7  D�  ��   ��  �       ��=       ���� �����  �  �         ����  F G          X$� �     n  ʊ  �   ��  �	       ��=       ���� #K  �  �  �         ����  2 3          �� �� x     �  }  �      �        ��>        ���� � �����  �  �         ����  4 5          �� �� y     �  �~  l�       �       ��>        ���� � �����  �  �         ����  6 7          �� �� z     �   �  �   ��  �       ��>        ���� � �����  �  �         ����  8 9          �� �� {     &  ��     ��  �       ��>       ���� � �����  �  �         ����  : ;          �� �� |     ]  ,�  h,   ��  �       ��>       ����  �����  �  �         ����  < =          �� �� }     �  ��  �A   ��  �       ��>       ���� �����  �  �         ����  ? @          �� �� ~     �  8�  W   ��  �       ��>       ���� �����  �  �         ����  A B          �� ��        ��  dl   ��  �       ��>       ���� �����  �  �         ����  C D          �� �� �     7  D�  ��   ��  �       ��>       ���� �����  �  �         ����  E F          �� �� �     n  ʊ  �   ��  �	       ��>       ���� #K  �  �  �         ����  & '          � �� x     �  }  �      �        ��?        ���� � �����  �  �         ����  ( )          � �� y     �  �~  l�       �       ��?        ���� � �����  �  �         ����  * +          � %�� z     �   �  �   ��  �       ��?        ���� � �����  �  �         ����  , -          � +�� {     &  ��     ��  �       ��?       ���� � �����  �  �         ����  . /          � 1 � |     ]  ,�  h,   ��  �       ��?       ����  �����  �  �         ����  0 1          � 7� }     �  ��  �A   ��  �       ��?       ���� �����  �  �         ����  2 3          � =� ~     �  8�  W   ��  �       ��?       ���� �����  �  �         ����  4 5          � C�        ��  dl   ��  �       ��?       ���� �����  �  �         ����  6 7          � I � �     7  D�  ��   ��  �       ��?       ���� �����  �  �         ����  8 9          � O(� �     n  ʊ  �   ��  �	       ��?       ���� #K  �  �  �         ����  5 6          hx� � x     �  }  �              ��@        ���� � �����  �  �         ����  7 8          o� � y     �  �~  l�              ��@        ���� � �����  �  �         ����  9 :          v�� � z     �   �  �   ��         ��@        ���� � �����  �  �         ����  ; <          }�� � {     &  ��     ��         ��@       ���� � �����  �  �         ����  = >          ��� � |     ]  ,�  h,   ��         ��@       ����  �����  �  �         ����  ? @          ��� � }     �  ��  �A   ��         ��@       ���� �����  �  �         ����  B C          ��� � ~     �  8�  W   ��         ��@       ���� �����  �  �         ����  D E          ��� �        ��  dl   ��         ��@       ���� �����  �  �         ����  F G          ��� � �     7  D�  ��   ��         ��@       ���� �����  �  �         ����  H I          ��� � �     n  ʊ  �   ��  	       ��@       ���� #K  �  �  �         ����  @ A          �� � x     J  �{  8�      .        ��A        ���� � �����  �  �         ����  B C          �� � y     �  
}  ��       .       ��A        ���� � �����  �  �         ����  D E          �$� � z     �  �~  ��   ��  .       ��A        ���� � �����  �  �         ����  G H          �*� � {     �  �  4   ��  .       ��A       ���� � �����  �  �         ����  I J          �0� � |     %  ��  �   ��  .       ��A       ����  �����  �  �         ����  K L          �6� � }     [  "�  �+   ��  .       ��A       ���� �����  �  �         ����  M N          �<� � ~     �  ��  0A   ��  .       ��A       ���� �����  �  �         ����  O P          B� �      �  .�  �V   ��  .       ��A       ���� �����  �  �         ����  R S          	H� � �     �  ��  �k   ��  .       ��A       ���� �����  �  �         ����  T U          N� � �     6  :�  ,�   ��  .	       ��A       ���� #K  �  �  �         ����  2 3          � �� x     J  �{  8�      ?        ��B        ���� � �����  �  �         ����  4 5          � �� y     �  
}  ��       ?       ��B        ���� � �����  �  �         ����  6 7          � �� z     �  �~  ��   ��  ?       ��B        ���� � �����  �  �         ����  8 9          � �� {     �  �  4   ��  ?       ��B       ���� � �����  �  �         ����  : ;          �  �� |     %  ��  �   ��  ?       ��B       ����  �����  �  �         ����  < =          � &�� }     [  "�  �+   ��  ?       ��B       ���� �����  �  �         ����  ? @          � ,�� ~     �  ��  0A   ��  ?       ��B       ���� �����  �  �         ����  A B          � 2��      �  .�  �V   ��  ?       ��B       ���� �����  �  �         ����  C D          � 8� �     �  ��  �k   ��  ?       ��B       ���� �����  �  �         ����  E F          � >
� �     6  :�  ,�   ��  ?	       ��B       ���� #K  �  �  �         ����  1 2          w� w� x     J  �{  8�      P        ��C        ���� � �����  �  �         ����  3 4          ~� ~� y     �  
}  ��       P       ��C        ���� � �����  �  �         ����  5 6          �� �� z     �  �~  ��   ��  P       ��C        ���� � �����  �  �         ����  7 8          �� �� {     �  �  4   ��  P       ��C       ���� � �����  �  �         ����  9 :          �� �� |     %  ��  �   ��  P       ��C       ����  �����  �  �         ����  ; <          �� �� }     [  "�  �+   ��  P       ��C       ���� �����  �  �         ����  > ?          �� �� ~     �  ��  0A   ��  P       ��C       ���� �����  �  �         ����  @ A          �� ��      �  .�  �V   ��  P       ��C       ���� �����  �  �         ����  B C          �� �� �     �  ��  �k   ��  P       ��C       ���� �����  �  �         ����  D E          �� �� �     6  :�  ,�   ��  P	       ��C       ���� #K  �  �  �         ����  % &          � �� x     J  �{  8�      a        ��D        ���� � �����  �  �         ����  ' (          � �� y     �  
}  ��       a       ��D        ���� � �����  �  �         ����  ) *          � �� z     �  �~  ��   ��  a       ��D        ���� � �����  �  �         ����  + ,          � "�� {     �  �  4   ��  a       ��D       ���� � �����  �  �         ����  - .          � (�� |     %  ��  �   ��  a       ��D       ����  �����  �  �         ����  / 0          � .�� }     [  "�  �+   ��  a       ��D       ���� �����  �  �         ����  1 2          � 4� ~     �  ��  0A   ��  a       ��D       ���� �����  �  �         ����  3 4          � :�      �  .�  �V   ��  a       ��D       ���� �����  �  �         ����  5 6          � @� �     �  ��  �k   ��  a       ��D       ���� �����  �  �         ����  7 8          � F� �     6  :�  ,�   ��  a	       ��D       ���� #K  �  �  �         ����  4 5          he� � x     J  �{  8�      r        ��E        ���� � �����  �  �         ����  6 7          ol� � y     �  
}  ��       r       ��E        ���� � �����  �  �         ����  8 9          vs� � z     �  �~  ��   ��  r       ��E        ���� � �����  �  �         ����  : ;          }z� � {     �  �  4   ��  r       ��E       ���� � �����  �  �         ����  < =          ��� � |     %  ��  �   ��  r       ��E       ����  �����  �  �         ����  > ?          ��� � }     [  "�  �+   ��  r       ��E       ���� �����  �  �         ����  A B          ��� � ~     �  ��  0A   ��  r       ��E       ���� �����  �  �         ����  C D          ��� �      �  .�  �V   ��  r       ��E       ���� �����  �  �         ����  E F          ��� � �     �  ��  �k   ��  r       ��E       ���� �����  �  �         ����  G H          ��� � �     6  :�  ,�   ��  r	       ��E       ���� #K  �  �  �         ����  A B          �� � x     �  4�  �      �      �   F        ���� � �����  �  �         ����  C D          �� � y     )  ��  ,       �     �   F        ���� � �����  �  �         ����  E F          �$� � z     `  @�  �-   ��  �     �   F        ���� � �����  �  �         ����  H I          �*� � {     �  Ƅ  �B   ��  �     �   F       ���� � �����  �  �         ����  J K          �0� � |     �  L�  (X   ��  �     �   F       ����  �����  �  �         ����  L M          6� � }       ҇  |m   ��  �     �   F       ���� �����  �  �         ����  N O          <� � ~     :  X�  Ђ   ��  �     �   F       ���� �����  �  �         ����  P Q          B� �      q  ފ  $�   ��  �     �   F       ���� �����  �  �         ����  S T          H� � �     �  d�  x�   ��  �     �   F       ���� �����  �  �         ����  U V          #N� � �     �  �  ��   ��  �	     �   F       ���� #K  �  �  �         ����  3 4          � �� x     �  4�  �      �      �   G        ���� � �����  �  �         ����  5 6          �  �� y     )  ��  ,       �     �   G        ���� � �����  �  �         ����  7 8          � &�� z     `  @�  �-   ��  �     �   G        ���� � �����  �  �         ����  9 :          � ,�� {     �  Ƅ  �B   ��  �     �   G       ���� � �����  �  �         ����  ; <          � 2�� |     �  L�  (X   ��  �     �   G       ����  �����  �  �         ����  = >          � 8�� }       ҇  |m   ��  �     �   G       ���� �����  �  �         ����  @ A          � >� ~     :  X�  Ђ   ��  �     �   G       ���� �����  �  �         ����  B C          � D�      q  ފ  $�   ��  �     �   G       ���� �����  �  �         ����  D E          � J� �     �  d�  x�   ��  �     �   G       ���� �����  �  �         ����  F G          � P� �     �  �  ��   ��  �	     �   G       ���� #K  �  �  �         ����  2 3          �� �� x     �  4�  �      �      �   H        ���� � �����  �  �         ����  4 5          �� �� y     )  ��  ,       �     �   H        ���� � �����  �  �         ����  6 7          �� �� z     `  @�  �-   ��  �     �   H        ���� � �����  �  �         ����  8 9          �� �� {     �  Ƅ  �B   ��  �     �   H       ���� � �����  �  �         ����  : ;          �� �� |     �  L�  (X   ��  �     �   H       ����  �����  �  �         ����  < =          �� �� }       ҇  |m   ��  �     �   H       ���� �����  �  �         ����  ? @          �� �� ~     :  X�  Ђ   ��  �     �   H       ���� �����  �  �         ����  A B          �� ��      q  ފ  $�   ��  �     �   H       ���� �����  �  �         ����  C D          �� �� �     �  d�  x�   ��  �     �   H       ���� �����  �  �         ����  E F          �� �� �     �  �  ��   ��  �	     �   H       ���� #K  �  �  �         ����  ' (          � � �� x     �  4�  �      �      �   I        ���� � �����  �  �         ����  ) *          � �� y     )  ��  ,       �     �   I        ���� � �����  �  �         ����  + ,          � 	�� z     `  @�  �-   ��  �     �   I        ���� � �����  �  �         ����  - .          � �� {     �  Ƅ  �B   ��  �     �   I       ���� � �����  �  �         ����  / 0          � �� |     �  L�  (X   ��  �     �   I       ����  �����  �  �         ����  1 2          � �� }       ҇  |m   ��  �     �   I       ���� �����  �  �         ����  3 4          � !�� ~     :  X�  Ђ   ��  �     �   I       ���� �����  �  �         ����  5 6          � '��      q  ފ  $�   ��  �     �   I       ���� �����  �  �         ����  7 8          � -�� �     �  d�  x�   ��  �     �   I       ���� �����  �  �         ����  9 :          � 3� �     �  �  ��   ��  �	     �   I       ���� #K  �  �  �         ����	  ? @           �� � x     �����  xD      �      �� ��J        ���� � �����  �  �         ����	  A B           �� � y     ����j�  �Y       �     �� ��J        ���� � �����  �  �         ����	  C D           �$� � z     ������   o   ��  �     �� ��J        ���� � �����  �  �         ����	  F G           �*� � {     ����v�  t�   ��  �     �� ��J       ���� � �����  �  �         ����	  H I           �0� � |     ������  ș   ��  �     �� ��J       ����  �����  �  �         ����	  J K           �6� � }     ������  �   ��  �     �� ��J       ���� �����  �  �         ����	  L M           �<� � ~     �����  p�   ��  �     �� ��J       ���� �����  �  �         ����	  N O           �B� �      ������  ��   ��  �     �� ��J       ���� �����  �  �         ����	  Q R           H� � �     �����  �   ��  �     �� ��J       ���� �����  �  �         ����	  S T           N� � �     ������  l   ��  �	     �� ��J       ���� #�����  �  �         ����	  2 3           � �� x     �����  xD      �      �� ��J        ���� � �����  �  �         ����	  4 5           � 	�� y     ����j�  �Y       �     �� ��J        ���� � �����  �  �         ����	  6 7           � �� z     ������   o   ��  �     �� ��J        ���� � �����  �  �         ����	  8 9           � �� {     ����v�  t�   ��  �     �� ��J       ���� � �����  �  �         ����	  : ;           � �� |     ������  ș   ��  �     �� ��J       ����  �����  �  �         ����	  < =           � !�� }     ������  �   ��  �     �� ��J       ���� �����  �  �         ����	  ? @           � '�� ~     �����  p�   ��  �     �� ��J       ���� �����  �  �         ����	  A B           � -��      ������  ��   ��  �     �� ��J       ���� �����  �  �         ����	  C D           � 3�� �     �����  �   ��  �     �� ��J       ���� �����  �  �         ����	  E F           � 9� �     ������  l   ��  �	     �� ��J       ���� #�����  �  �         ����	  1 2           r� r� x     �����  xD            �� ��J        ���� � �����  �  �         ����	  3 4           y� y� y     ����j�  �Y            �� ��J        ���� � �����  �  �         ����	  5 6           �� �� z     ������   o   ��       �� ��J        ���� � �����  �  �         ����	  7 8           �� �� {     ����v�  t�   ��       �� ��J       ���� � �����  �  �         ����	  9 :           �� �� |     ������  ș   ��       �� ��J       ����  �����  �  �         ����	  ; <           �� �� }     ������  �   ��       �� ��J       ���� �����  �  �         ����	  > ?           �� �� ~     �����  p�   ��       �� ��J       ���� �����  �  �         ����	  @ A           �� ��      ������  ��   ��       �� ��J       ���� �����  �  �         ����	  B C           �� �� �     �����  �   ��       �� ��J       ���� �����  �  �         ����	  D E           �� �� �     ������  l   ��  	     �� ��J       ���� #�����  �  �         ����	  & '           � � �� x     �����  xD            �� ��J        ���� � �����  �  �         ����	  ( )           �  �� y     ����j�  �Y            �� ��J        ���� � �����  �  �         ����	  * +           � �� z     ������   o   ��       �� ��J        ���� � �����  �  �         ����	  , -           � �� {     ����v�  t�   ��       �� ��J       ���� � �����  �  �         ����	  . /           � �� |     ������  ș   ��       �� ��J       ����  �����  �  �         ����	  0 1           � �� }     ������  �   ��       �� ��J       ���� �����  �  �         ����	  2 3           � �� ~     �����  p�   ��       �� ��J       ���� �����  �  �         ����	  4 5           � $��      ������  ��   ��       �� ��J       ���� �����  �  �         ����	  6 7           � *�� �     �����  �   ��       �� ��J       ���� �����  �  �         ����	  8 9           � 0� �     ������  l   ��  	     �� ��J       ���� #�����  �  �         ����	  3 4           he� � x     �����  xD      %      ��  ��J        ���� � �����  �  �         ����	  5 6           ol� � y     ����j�  �Y       %     ��  ��J        ���� � �����  �  �         ����	  7 8           vs� � z     ������   o   ��  %     ��  ��J        ���� � �����  �  �         ����	  9 :           }z� � {     ����v�  t�   ��  %     ��  ��J       ���� � �����  �  �         ����	  ; <           ��� � |     ������  ș   ��  %     ��  ��J       ����  �����  �  �         ����	  = >           ��� � }     ������  �   ��  %     ��  ��J       ���� �����  �  �         ����	  @ A           ��� � ~     �����  p�   ��  %     ��  ��J       ���� �����  �  �         ����	  B C           ��� �      ������  ��   ��  %     ��  ��J       ���� �����  �  �         ����	  D E           ��� � �     �����  �   ��  %     ��  ��J       ���� �����  �  �         ����	  F G           ��� � �     ������  l   ��  %	     ��  ��J       ���� #�����  �  �         ����
  @ A           �� � x     ����T�  �.      C      �� ��K        ���� � �����  �  �         ����
  B C           �� � y     ����ڄ  �C       C     �� ��K        ���� � �����  �  �         ����
  D E           �$� � z     ����`�  @Y   ��  C     �� ��K        ���� � �����  �  �         ����
  G H           �*� � {     �����  �n   ��  C     �� ��K       ���� � �����  �  �         ����
  I J           �0� � |     ����l�  �   ��  C     �� ��K       ����  �����  �  �         ����
  K L           �6� � }     �����  <�   ��  C     �� ��K       ���� �����  �  �         ����
  M N           <� � ~     ����x�  ��   ��  C     �� ��K       ���� �����  �  �         ����
  O P           	B� �      ������  ��   ��  C     �� ��K       ���� �����  �  �         ����
  R S           H� � �     ������  8�   ��  C     �� ��K       ���� �����  �  �         ����
  T U           N� � �     ����
�  ��   ��  C	     �� ��K       ���� #�����  �  �         ����
  2 3           � �� x     ����T�  �.      R      �� ��K        ���� � �����  �  �         ����
  4 5           � �� y     ����ڄ  �C       R     �� ��K        ���� � �����  �  �         ����
  6 7           � �� z     ����`�  @Y   ��  R     �� ��K        ���� � �����  �  �         ����
  8 9           � "�� {     �����  �n   ��  R     �� ��K       ���� � �����  �  �         ����
  : ;           � (�� |     ����l�  �   ��  R     �� ��K       ����  �����  �  �         ����
  < =           � .�� }     �����  <�   ��  R     �� ��K       ���� �����  �  �         ����
  ? @           � 4�� ~     ����x�  ��   ��  R     �� ��K       ���� �����  �  �         ����
  A B           � :�      ������  ��   ��  R     �� ��K       ���� �����  �  �         ����
  C D           � @
� �     ������  8�   ��  R     �� ��K       ���� �����  �  �         ����
  E F           � F� �     ����
�  ��   ��  R	     �� ��K       ���� #�����  �  �         ����
  1 2           � � x     ����T�  �.      a      �� ��K        ���� � �����  �  �         ����
  3 4           �� �� y     ����ڄ  �C       a     �� ��K        ���� � �����  �  �         ����
  5 6           �� �� z     ����`�  @Y   ��  a     �� ��K        ���� � �����  �  �         ����
  7 8           �� �� {     �����  �n   ��  a     �� ��K       ���� � �����  �  �         ����
  9 :           �� �� |     ����l�  �   ��  a     �� ��K       ����  �����  �  �         ����
  ; <           �� �� }     �����  <�   ��  a     �� ��K       ���� �����  �  �         ����
  > ?           �� �� ~     ����x�  ��   ��  a     �� ��K       ���� �����  �  �         ����
  @ A           �� ��      ������  ��   ��  a     �� ��K       ���� �����  �  �         ����
  B C           �� �� �     ������  8�   ��  a     �� ��K       ���� �����  �  �         ����
  D E           �� �� �     ����
�  ��   ��  a	     �� ��K       ���� #�����  �  �         ����
  & '           � �� x     ����T�  �.      p      �� ��K        ���� � �����  �  �         ����
  ( )           � 	�� y     ����ڄ  �C       p     �� ��K        ���� � �����  �  �         ����
  * +           � �� z     ����`�  @Y   ��  p     �� ��K        ���� � �����  �  �         ����
  , -           � �� {     �����  �n   ��  p     �� ��K       ���� � �����  �  �         ����
  . /           � �� |     ����l�  �   ��  p     �� ��K       ����  �����  �  �         ����
  0 1           � !�� }     �����  <�   ��  p     �� ��K       ���� �����  �  �         ����
  2 3           � '�� ~     ����x�  ��   ��  p     �� ��K       ���� �����  �  �         ����
  4 5           � -��      ������  ��   ��  p     �� ��K       ���� �����  �  �         ����
  6 7           � 3� �     ������  8�   ��  p     �� ��K       ���� �����  �  �         ����
  8 9           � 9� �     ����
�  ��   ��  p	     �� ��K       ���� #�����  �  �         ����
  4 5           hm� � x     ����T�  �.            ��  ��K        ���� � �����  �  �         ����
  6 7           ot� � y     ����ڄ  �C            ��  ��K        ���� � �����  �  �         ����
  8 9           v{� � z     ����`�  @Y   ��       ��  ��K        ���� � �����  �  �         ����
  : ;           }�� � {     �����  �n   ��       ��  ��K       ���� � �����  �  �         ����
  < =           ��� � |     ����l�  �   ��       ��  ��K       ����  �����  �  �         ����
  > ?           ��� � }     �����  <�   ��       ��  ��K       ���� �����  �  �         ����
  A B           ��� � ~     ����x�  ��   ��       ��  ��K       ���� �����  �  �         ����
  C D           ��� �      ������  ��   ��       ��  ��K       ���� �����  �  �         ����
  E F           ��� � �     ������  8�   ��       ��  ��K       ���� �����  �  �         ����
  G H           ��� � �     ����
�  ��   ��  	     ��  ��K       ���� #�����  �  �         ����  A B           �� � x     �����x  �      �      �� ��L        ���� � �����  �  �         ����  C D           �� � y     ����Nz  D�       �     �� ��L        ���� � �����  �  �         ����  E F           �$� � z     �����{  ��   ��  �     �� ��L        ���� � �����  �  �         ����  H I           �*� � {     ����Z}  ��   ��  �     �� ��L       ���� � �����  �  �         ����  J K           �0� � |     �����~  @�   ��  �     �� ��L       ����  �����  �  �         ����  L M           6� � }     ����f�  �   ��  �     �� ��L       ���� �����  �  �         ����  N O           <� � ~     �����  �   ��  �     �� ��L       ���� �����  �  �         ����  P Q           B� �      ����r�  <0   ��  �     �� ��L       ���� �����  �  �         ����  S T           H� � �     ������  �E   ��  �     �� ��L       ���� �����  �  �         ����  U V           &N� � �     ����~�  �Z   ��  �	     �� ��L       ���� #�����  �  �         ����  3 4           � �� x     �����x  �      �      �� ��L        ���� � �����  �  �         ����  5 6           � #�� y     ����Nz  D�       �     �� ��L        ���� � �����  �  �         ����  7 8           � )�� z     �����{  ��   ��  �     �� ��L        ���� � �����  �  �         ����  9 :           � /�� {     ����Z}  ��   ��  �     �� ��L       ���� � �����  �  �         ����  ; <           � 5�� |     �����~  @�   ��  �     �� ��L       ����  �����  �  �         ����  = >           � ;�� }     ����f�  �   ��  �     �� ��L       ���� �����  �  �         ����  @ A           � A� ~     �����  �   ��  �     �� ��L       ���� �����  �  �         ����  B C           � G�      ����r�  <0   ��  �     �� ��L       ���� �����  �  �         ����  D E           � M� �     ������  �E   ��  �     �� ��L       ���� �����  �  �         ����  F G           S� �     ����~�  �Z   ��  �	     �� ��L       ���� #�����  �  �         ����  2 3           �� �� x     �����x  �      �      �� ��L        ���� � �����  �  �         ����  4 5           �� �� y     ����Nz  D�       �     �� ��L        ���� � �����  �  �         ����  6 7           �� �� z     �����{  ��   ��  �     �� ��L        ���� � �����  �  �         ����  8 9           �� �� {     ����Z}  ��   ��  �     �� ��L       ���� � �����  �  �         ����  : ;           �� �� |     �����~  @�   ��  �     �� ��L       ����  �����  �  �         ����  < =           �� �� }     ����f�  �   ��  �     �� ��L       ���� �����  �  �         ����  ? @           �� �� ~     �����  �   ��  �     �� ��L       ���� �����  �  �         ����  A B           �� ��      ����r�  <0   ��  �     �� ��L       ���� �����  �  �         ����  C D           �� �� �     ������  �E   ��  �     �� ��L       ���� �����  �  �         ����  E F           �� �� �     ����~�  �Z   ��  �	     �� ��L       ���� #�����  �  �         ����  & '           � �� x     �����x  �      �      �� ��L        ���� � �����  �  �         ����  ( )           � �� y     ����Nz  D�       �     �� ��L        ���� � �����  �  �         ����  * +           � �� z     �����{  ��   ��  �     �� ��L        ���� � �����  �  �         ����  , -           � �� {     ����Z}  ��   ��  �     �� ��L       ���� � �����  �  �         ����  . /           � $�� |     �����~  @�   ��  �     �� ��L       ����  �����  �  �         ����  0 1           � *�� }     ����f�  �   ��  �     �� ��L       ���� �����  �  �         ����  2 3           � 0�� ~     �����  �   ��  �     �� ��L       ���� �����  �  �         ����  4 5           � 6�      ����r�  <0   ��  �     �� ��L       ���� �����  �  �         ����  6 7           � <� �     ������  �E   ��  �     �� ��L       ���� �����  �  �         ����  8 9           � B� �     ����~�  �Z   ��  �	     �� ��L       ���� #�����  �  �         ����  5 6           hu� � x     �����x  �      �      ��  ��L        ���� � �����  �  �         ����  7 8           o|� � y     ����Nz  D�       �     ��  ��L        ���� � �����  �  �         ����  9 :           v�� � z     �����{  ��   ��  �     ��  ��L        ���� � �����  �  �         ����  ; <           }�� � {     ����Z}  ��   ��  �     ��  ��L       ���� � �����  �  �         ����  = >           ��� � |     �����~  @�   ��  �     ��  ��L       ����  �����  �  �         ����  ? @           ��� � }     ����f�  �   ��  �     ��  ��L       ���� �����  �  �         ����  B C           ��� � ~     �����  �   ��  �     ��  ��L       ���� �����  �  �         ����  D E           ��� �      ����r�  <0   ��  �     ��  ��L       ���� �����  �  �         ����  F G           ��� � �     ������  �E   ��  �     ��  ��L       ���� �����  �  �         ����  H I           ��� � �     ����~�  �Z   ��  �	     ��  ��L       ���� #�����  �  �         ����  B C           �� � x     ����t�  XZ      �      �� ��M        ���� � �����  �  �         ����  D E           �� � y     ������  �o       �     �� ��M        ���� � �����  �  �         ����  F G           �$� � z     ������   �   ��  �     �� ��M        ���� � �����  �  �         ����  I J           *� � {     �����  T�   ��  �     �� ��M       ���� � �����  �  �         ����  K L           0� � |     ������  ��   ��  �     �� ��M       ����  �����  �  �         ����  M N           6� � }     �����  ��   ��  �     �� ��M       ���� �����  �  �         ����  O P           <� � ~     ������  P�   ��  �     �� ��M       ���� �����  �  �         ����  Q R           #B� �      �����  ��   ��  �     �� ��M       ���� �����  �  �         ����  T U           +H� � �     ������  �   ��  �     �� ��M       ���� �����  �  �         ����  V W           3N� � �     ����*�  L   ��  �	     �� ��M       ���� #�����  �  �         ����  3 4           � *�� x     ����t�  XZ            �� ��M        ���� � �����  �  �         ����  5 6           � 0�� y     ������  �o            �� ��M        ���� � �����  �  �         ����  7 8           � 6�� z     ������   �   ��       �� ��M        ���� � �����  �  �         ����  9 :           � <�� {     �����  T�   ��       �� ��M       ���� � �����  �  �         ����  ; <           � B� |     ������  ��   ��       �� ��M       ����  �����  �  �         ����  = >           � H� }     �����  ��   ��       �� ��M       ���� �����  �  �         ����  @ A           � N� ~     ������  P�   ��       �� ��M       ���� �����  �  �         ����  B C           T�      �����  ��   ��       �� ��M       ���� �����  �  �         ����  D E           	Z$� �     ������  �   ��       �� ��M       ���� �����  �  �         ����  F G           `,� �     ����*�  L   ��  	     �� ��M       ���� #�����  �  �         ����  2 3           �� �� x     ����t�  XZ            �� ��M        ���� � �����  �  �         ����  4 5           �� �� y     ������  �o            �� ��M        ���� � �����  �  �         ����  6 7           �� �� z     ������   �   ��       �� ��M        ���� � �����  �  �         ����  8 9           �� �� {     �����  T�   ��       �� ��M       ���� � �����  �  �         ����  : ;           �� �� |     ������  ��   ��       �� ��M       ����  �����  �  �         ����  < =           �� �� }     �����  ��   ��       �� ��M       ���� �����  �  �         ����  ? @           �� �� ~     ������  P�   ��       �� ��M       ���� �����  �  �         ����  A B           �� ��      �����  ��   ��       �� ��M       ���� �����  �  �         ����  C D           �� �� �     ������  �   ��       �� ��M       ���� �����  �  �         ����  E F           �� �� �     ����*�  L   ��  	     �� ��M       ���� #�����  �  �         ����  & '           � �� x     ����t�  XZ      $      �� ��M        ���� � �����  �  �         ����  ( )           � �� y     ������  �o       $     �� ��M        ���� � �����  �  �         ����  * +           � !�� z     ������   �   ��  $     �� ��M        ���� � �����  �  �         ����  , -           � '�� {     �����  T�   ��  $     �� ��M       ���� � �����  �  �         ����  . /           � -�� |     ������  ��   ��  $     �� ��M       ����  �����  �  �         ����  0 1           � 3�� }     �����  ��   ��  $     �� ��M       ���� �����  �  �         ����  2 3           � 9� ~     ������  P�   ��  $     �� ��M       ���� �����  �  �         ����  4 5           � ?�      �����  ��   ��  $     �� ��M       ���� �����  �  �         ����  6 7           � E� �     ������  �   ��  $     �� ��M       ���� �����  �  �         ����  8 9           � K� �     ����*�  L   ��  $	     �� ��M       ���� #�����  �  �         ����  5 6           h}� � x     ����t�  XZ      3      ��  ��M        ���� � �����  �  �         ����  7 8           o�� � y     ������  �o       3     ��  ��M        ���� � �����  �  �         ����  9 :           v�� � z     ������   �   ��  3     ��  ��M        ���� � �����  �  �         ����  ; <           }�� � {     �����  T�   ��  3     ��  ��M       ���� � �����  �  �         ����  = >           ��� � |     ������  ��   ��  3     ��  ��M       ����  �����  �  �         ����  ? @           ��� � }     �����  ��   ��  3     ��  ��M       ���� �����  �  �         ����  B C           ��� � ~     ������  P�   ��  3     ��  ��M       ���� �����  �  �         ����  D E           ��� �      �����  ��   ��  3     ��  ��M       ���� �����  �  �         ����  F G           ��� � �     ������  �   ��  3     ��  ��M       ���� �����  �  �         ����  H I           ��� � �     ����*�  L   ��  3	     ��  ��M       ���� #�����  �  �         ����  B C           �� � x     �����  8p      Q      �� ��N        ���� � �����  �  �         ����  D E           �� � y     ������  ��       Q     �� ��N        ���� � �����  �  �         ����  F G           �$� � z     �����  ��   ��  Q     �� ��N        ���� � �����  �  �         ����  I J           *� � {     ������  4�   ��  Q     �� ��N       ���� � �����  �  �         ����  K L           0� � |     �����  ��   ��  Q     �� ��N       ����  �����  �  �         ����  M N           6� � }     ������  ��   ��  Q     �� ��N       ���� �����  �  �         ����  O P           <� � ~     ����(�  0�   ��  Q     �� ��N       ���� �����  �  �         ����  Q R           &B� �      ������  �   ��  Q     �� ��N       ���� �����  �  �         ����  T U           .H� � �     ����4�  �   ��  Q     �� ��N       ���� �����  �  �         ����  V W           6N� � �     ������  ,0   ��  Q	     �� ��N       ���� #�����  �  �         ����  3 4           � -�� x     �����  8p      `      �� ��N        ���� � �����  �  �         ����  5 6           � 3�� y     ������  ��       `     �� ��N        ���� � �����  �  �         ����  7 8           � 9�� z     �����  ��   ��  `     �� ��N        ���� � �����  �  �         ����  9 :           � ?�� {     ������  4�   ��  `     �� ��N       ���� � �����  �  �         ����  ; <           � E� |     �����  ��   ��  `     �� ��N       ����  �����  �  �         ����  = >           � K� }     ������  ��   ��  `     �� ��N       ���� �����  �  �         ����  @ A           Q� ~     ����(�  0�   ��  `     �� ��N       ���� �����  �  �         ����  B C           W�      ������  �   ��  `     �� ��N       ���� �����  �  �         ����  D E           ]'� �     ����4�  �   ��  `     �� ��N       ���� �����  �  �         ����  F G           c/� �     ������  ,0   ��  `	     �� ��N       ���� #�����  �  �         ����  2 3           �� �� x     �����  8p      o      �� ��N        ���� � �����  �            ����  4 5           �� �� y     ������  ��       o     �� ��N        ���� � �����  �            ����  6 7           �� �� z     �����  ��   ��  o     �� ��N        ���� � �����  �            ����  8 9           �� �� {     ������  4�   ��  o     �� ��N       ���� � �����  �            ����  : ;           �� �� |     �����  ��   ��  o     �� ��N       ����  �����  �            ����  < =           �� �� }     ������  ��   ��  o     �� ��N       ���� �����  �            ����  ? @           �� �� ~     ����(�  0�   ��  o     �� ��N       ���� �����  �            ����  A B           �� ��      ������  �   ��  o     �� ��N       ���� �����  �            ����  C D           �� �� �     ����4�  �   ��  o     �� ��N       ���� �����  �            ����  E F           �� �� �     ������  ,0   ��  o	     �� ��N       ���� #�����  �            ����  & '           � �� x     �����  8p      ~      �� ��N        ���� � �����  �           ����  ( )           � �� y     ������  ��       ~     �� ��N        ���� � �����  �           ����  * +           � $�� z     �����  ��   ��  ~     �� ��N        ���� � �����  �           ����  , -           � *�� {     ������  4�   ��  ~     �� ��N       ���� � �����  �           ����  . /           � 0�� |     �����  ��   ��  ~     �� ��N       ����  �����  �           ����  0 1           � 6� }     ������  ��   ��  ~     �� ��N       ���� �����  �           ����  2 3           � <
� ~     ����(�  0�   ��  ~     �� ��N       ���� �����  �           ����  4 5           � B�      ������  �   ��  ~     �� ��N       ���� �����  �           ����  6 7           � H� �     ����4�  �   ��  ~     �� ��N       ���� �����  �           ����  8 9           N"� �     ������  ,0   ��  ~	     �� ��N       ���� #�����  �           ����  5 6           h� � x     �����  8p      �      ��  ��N        ���� � �����  �           ����  7 8           o�� � y     ������  ��       �     ��  ��N        ���� � �����  �           ����  9 :           v�� � z     �����  ��   ��  �     ��  ��N        ���� � �����  �           ����  ; <           }�� � {     ������  4�   ��  �     ��  ��N       ���� � �����  �           ����  = >           ��� � |     �����  ��   ��  �     ��  ��N       ����  �����  �           ����  ? @           ��� � }     ������  ��   ��  �     ��  ��N       ���� �����  �           ����  B C           ��� � ~     ����(�  0�   ��  �     ��  ��N       ���� �����  �           ����  D E           ��� �      ������  �   ��  �     ��  ��N       ���� �����  �           ����  F G           ��� � �     ����4�  �   ��  �     ��  ��N       ���� �����  �           ����  H I           ��� � �     ������  ,0   ��  �	     ��  ��N       ���� #�����  �            s g                ��O�n     ������  %�       �      ��$ ���         ����   ����������������        t g                �i�}     ����h�  �       �      ��$ ���         ����   ����������������        u g                �C>n     ������  %�       �      ��% ���         ����   ����������������        v g                �a?Z}     ����h�  �       �      ��% ���         ����   ����������������        w g                ���n     ������  %�             ��& ��        ����   ����������������        x g                -���}     ����h�  �       	      ��& ��        ����   ����������������        y g                �%.An     ������  %�       !      ��' ���        ����   ����������������        z g                �J`T}     ����h�  �       "      ��' ���        ����   ����������������        { g                ��cn     ������  %�       :      ��( ��        ����   ����������������        | g                ���~}     ����h�  �       ;      ��( ��        ����   ����������������       ����{ ��                            �� '  '        �      ��e ��O        ������  ����������������       ����| ��                            �����a  �a       �      �� ��P        ������  ����������������       ����z ��                            ����'  @�        �      ��f ��Q        ������  ����������������        ��t ��                           ����'   N       ^      �� ��R        ������  ����������������        ��y ���td                     �� @B @B      r      �� ��S        ������  ����������������        ��y ��t<x _  R               �� �O �O      s      �� ��S        ������  ����������������        ��y ��<� '  �               �" �\ �\      t      �� ��S        ������  ����������������        ��y ���� �  �                q  j  j      u      �� ��S        ������  ����������������        ��y ����� �  �                � @w @w      v      �� ��S        ������  ����������������        ��y ���hd �  �               �I `� `�      w      �� ��S        ������  ����������������        ��y ��0�n _ �               � �� ��      x      �� ��S        ������  ����������������        ��y ����x ' �               0� �� ��      y      �� ��S        ������  ����������������        ��y ��P� � �               P4            z      �� ��S        ������  ����������������        ��y ����� �                p� `# `#      {      �� ��S        ������  ����������������        ��y ����P ' �               @ �� ��      |      �� ��S        ������  ����������������        ��y ���hZ ' �               `[ ��! ��!      }      �� ��S        ������  ����������������        ��y ��h0d ' �               ��  �$  �$      ~      �� ��S        ������  ����������������        ��y ��0�n � �               �� @�' @�'            �� ��S        ������  ����������������        ��y ����x �                �E ��* ��*      �      �� ��S        ������  ����������������        ��y ��0�< � X               �� �%& �%&      �      �� ��S        ������  ����������������        ��y ����F � b               � �2) �2)      �      �� ��S        ������  ����������������        ��y ����P � l               �l  @,  @,      �      �� ��S        ������  ����������������        ��y ���PZ � v               � `M/ `M/      �      �� ��S        ������  ����������������        ��y ��Pd � �               	 �Z2 �Z2      �      �� ��S        ������  ����������������       ����� ��                            �����  �        G      ��g ��T        ������  ����������������       ����� ��                            �����  �        H      ��g ��T        ������  ����������������       ����� ��                            �����  �        I      ��g ��T        ������  ����������������       ����� ��                            �����  �        J      ��g ��T        ������  ����������������       ����� ��                            �����  �        K      ��g ��T        ������  ����������������        } g                    
       �����   �        <      ��) ��U        ����   ����������������        ~ g                            ����B  �        =      ��) ��U        ����   ����������������         g                 ( " .        ����[  l        >      ��) ��U        ����   ����������������        � g                 1 - = (       ����'  �#        ?      ��) ��U        ����   ����������������        � g                 < 9 M 3       �����
  �?        @      ��) ��U        ����   ����������������        � g                 G F ^ >       �����  �g        A      ��) ��U        ����   ����������������        � g                 T T p J       �����  �        B      ��) ��U        ����   ����������������        � g                 c c � W       ����U  ��        C      ��) ��U        ����   ����������������        � g                 r t � d       �����  @<       D      ��) ��U        ����	   ����������������        � g                 � � � �       �����?  }       E      ��) ��U        ����
   ����������������        � g                 � � � ~       ����O.  �+       F      ��) ��U        ����   ����������������        � g                 � � � �       �����6  �       G      ��) ��U        ����   ����������������        � g                 � � � q       �����&  ʨ       H      ��) ��U        ����   ����������������        � g                 � � �       �����I  �O       I      ��) ��U        ����   ����������������        � g                 � � �       ����T  A       J      ��) ��U        ����   ����������������        � g                 � 5�       ����A_  QS       K      ��) ��U        ����   ����������������        � g                 %W�       ����$k  ��       L      ��) ��U        ����   ����������������        � g                 *Fy�       �����w  ��       M      ��) ��U        ����   ����������������        � g                 Eg�      �����  <d
       N      ��) ��U        ����   ����������������        � g                 `��#      ������  �       O      ��) ��U        ����   ����������������        � g                 |��;      ������  ��       P      ��) ��U        ����   ����������������        � g                 ��,T      �����  p�       Q      ��) ��U        ����   ����������������        � g                 ��hn      ����%�  x       R      ��) ��U        ����   ����������������       �����                               ����
   '  ;     �      �� ��V        ������  ����������������        ����                 ) )         	      �       x        ��W        ���� � ������������          ����                 ) .            >  |       x       ��W        ���� � ������������          ����                 ) 3            \  �       x       ��W        ���� � ������������          ����     	            ) 8            z  �       x       ��W       ���� � ������������          ����    
             ) =            �  0       x       ��W       ���� � ������������          ����                 ) B            �  l       x       ��W       ���� � ������������          ����                 ) G            �  �       x       ��W       ���� � ������������          ����                 ) L            �  �       x       ��W       ���� � ������������          ����                 ) Q                      x       ��W       ���� � ������������          ����                 ) V            .  \       x	       ��W       ���� � ������������          ����                 $ D         #   �  �       y        ��X        ���� � ������������          ����     	            ' I         %   �  �       y       ��X        ���� � ������������          ����    
             * N         '     Z       y       ��X        ���� � ������������          ����                 - S         )   Z         y       ��X       ���� � ������������          ����                 0 X         *   �  �       y       ��X       ���� � ������������          ����                 3 ]         ,   �  v       y       ��X       ���� � ������������          ����                 6 b         .     *       y       ��X       ���� � ������������          ����                 9 g         0   J  �       y       ��X       ���� � ������������          ����                 < l         2   �  �       y       ��X       ���� � ������������          ����                 ? q         3   �  F       y	       ��X       ���� � ������������          ����    
            + ^         N   �  �       z        ��Y        ���� � ������������         ����               ! / c         R     0        z       ��Y        ���� � ������������         ����               $ 3 h         V   f  �!       z       ��Y        ���� � ������������         ����               ' 7 m         Y   �   #       z       ��Y       ���� � ������������         ����               * ; r         ]   	  h$       z       ��Y       ���� � ������������         ����               - ? w         `   t	  �%       z       ��Y       ���� � ������������         ����               0 C |         d   �	  8'       z       ��Y       ���� � ������������         ����               3 G �         h   (
  �(       z       ��Y       ���� � ������������         ����               6 K �         k   �
  *       z       ��Y       ���� � ������������         ����               9 O �         o   �
  p+       z	       ��Y       ���� � ������������          ����               & < w        �   D  T=       {        ��Z        ���� � ������������         ����               ) @ }        �   �  �?       {       ��Z        ���� � ������������         ����               , D �         �   4  B       {       ��Z        ���� � ������������         ����               / H � #       �   �  \D       {       ��Z       ���� � ������������         ����               2 L � &       �   $  �F       {       ��Z       ���� � ������������         ����               5 P � )       �   �  I       {       ��Z       ���� � ������������         ����               8 T � ,       �     dK       {       ��Z       ���� � ������������         ����               ; X � /       �   �  �M       {       ��Z       ���� � ������������         ����                > \ � 2       �     P       {       ��Z       ���� � ������������         ����    ! "          A ` � 5       �   |  lR       {	       ��Z       ���� � ������������          ����               - L � !         \  (n       |        ��[        ���� � ������������         ����               0 P � $       #  �  �q       |       ��[        ���� � ������������         ����               3 T � '       ,  �  0u       |       ��[        ���� � ������������         ����               6 X � *       5    �x       |       ��[       ���� � ������������         ����               9 \ � -       >  �  8|       |       ��[       ���� � ������������         ����               < ` � 0       G  J  �       |       ��[       ���� � ������������         ����                ? d � 3       P  �  @�       |       ��[       ���� � ������������         ����    ! "          B h � 6       Y  v  Ć       |       ��[       ���� � ������������         ����    # $          E l � 9       b    H�    
   |       ��[       ���� � ������������         ����    % &          H p � <       k  �  ̍    	   |	       ��[       ���� � ������������          ����               4 [ � (       �  �  ֵ       }        ��\        ���� � ������������         ����               8 _ � +       �  �  º       }       ��\        ���� � ������������         ����               < c � .       �  b  ��       }       ��\        ���� � ������������         ����               @ g � 1       �    ��       }       ��\       ���� � ������������         ����               D k � 4         �  ��       }       ��\       ���� � ������������         ����    ! "          H o � 7         ~  r�       }       ��\       ���� � ������������         ����    # $          L s � :         2  ^�       }       ��\       ���� � ������������         ����    % &          P w � =       )  �  J�    	   }       ��\       ���� � ������������         ����    ' (          T { � @       6  �  6�       }       ��\       ���� � ������������         ����    ) *          X  � C       B  N   "�       }	       ��\       ���� � ������������         ����               D j � .       �  #  �      ~        ��]        ���� � �����  �  	         ����               H o � 2       �  �#  �      ~       ��]        ���� � �����  �  	         ����               L t � 6       �  �$  &      ~       ��]        ���� � �����  �  	         ����      !          P y � :         �%  �,      ~       ��]       ���� � �����  �  	         ����    " #          T ~ � >         f&  03      ~       ��]       ���� � �����  �  	         ����    $ %          X � � B       #  8'  �9   	   ~       ��]       ���� � �����  �  	         ����    ' (          \ �  F       4  
(  P@      ~       ��]       ���� � �����  �  	         ����    ) *          ` � J       D  �(  �F      ~       ��]       ���� � �����  �  	         ����    + ,          d � N       U  �)  pM      ~       ��]       ���� � �����  �  	         ����    - .          h � R       f  �*   T      ~	       ��]       ���� � �����  �  	         ����               T � � >         �-  �              ��^        ���� � �����  �  
         ����      !          X � B       4  �.  x�             ��^        ���� � �����  �  
         ����    " #          \ � 
F       J  �/  �             ��^        ���� � �����  �  
         ����    $ %          ` � J       _  �0  X�   	          ��^       ���� � �����  �  
         ����    & '          d � N       u  �1  Ƚ             ��^       ���� � �����  �  
         ����    ( )          h � R       �  x2  8�             ��^       ���� � �����  �  
         ����    + ,          l � &V       �  h3  ��             ��^       ���� � �����  �  
         ����    - .          p � -Z       �  X4  �             ��^       ���� � �����  �  
         ����    / 0          t � 4^       �  H5  ��             ��^       ���� � �����  �  
         ����    1 2          x � ;b       �  86  ��      	       ��^       ���� � -  �  �  
         ����    " #          c � %M       �  �9  �C      �      	  ��_        ����	 � �����  �           ����    $ %          g � ,Q       �  ;  <N   
   �     	  ��_        ����	 � �����  �           ����    & '          k � 3U         <  �X      �     	  ��_        ����	 � �����  �           ����    ( )          o � :Y         "=  Tc      �     	  ��_       ����	 � �����  �           ����    * +          s � A]       8  0>  �m      �     	  ��_       ����	 � �����  �           ����    , -          w � Ha       S  >?  lx      �     	  ��_       ����	 � �����  �           ����    / 0          { � Oe       n  L@  ��      �     	  ��_       ����	 � �����  �           ����    1 2           � Vi       �  ZA  ��      �     	  ��_       ����	 � �����  �           ����    3 4          � � ]m       �  hB  �       �     	  ��_       ����	 � �����  �           ����    5 6          � � dq       �  vC  ��   ��  �	     	  ��_       ����	 � 7  �  �           ����    & '          r � M\       �  �G  z   	   �      
  ��`        ����
 � �����  �           ����    ( )          w � T`         �H  ^!      �     
  ��`        ����
 � �����  �           ����    * +          | � [d       $  J  B.      �     
  ��`        ����
 � �����  �           ����    , -          � � bh       E  2K  &;      �     
  ��`       ����
 � �����  �           ����    . /          � � il       f  ^L  
H      �     
  ��`       ����
 � �����  �           ����    0 1          � � pp       �  �M  �T      �     
  ��`       ����
 � �����  �           ����    3 4          � � wt       �  �N  �a      �     
  ��`       ����
 � �����  �           ����    5 6          � � ~x       �  �O  �n   ��  �     
  ��`       ����
 � �����  �           ����    7 8          � � �|       �  Q  �{   ��  �     
  ��`       ����
 � �����  �           ����    9 :          � � ��       	  :R  ~�   ��  �	     
  ��`       ����
 7  �  �           ����    * +          � � tj d     n
  �V  �      �        ��a        ���� � �����  �           ����    , -          � � {o e     �
  4X  p"      �       ��a        ���� � �����  �           ����    . /          � � �t f     �
  ~Y  �1      �       ��a        ���� � �����  �           ����    0 1          � � �y g     �
  �Z  `A      �       ��a       ���� � �����  �           ����    2 3          � � �~ h       \  �P      �       ��a       ���� � �����  �           ����    4 5          � � �� i     4  \]  P`   ��  �       ��a       ���� � �����  �           ����    7 8          � � �� j     [  �^  �o   ��  �       ��a       ���� � �����  �           ����    9 :          � � �� k     �  �_  @   ��  �       ��a       ���� � �����  �           ����    ; <          � � �� l     �  :a  ��   ��  �       ��a       ���� �����  �           ����    = >          � � �� m     �  �b  0�   ��  �	       ��a       ���� A  �  �           ����    . /          � � �� n     z  �g  �C      �        ��b        ���� � �����  �           ����    0 1          � � �� o     �  i  V      �       ��b        ���� � �����  �           ����    2 3          � � �� p     �  |j  Lh      �       ��b        ���� � �����  �           ����    4 5          � � �� q       �k  �z   ��  �       ��b       ���� � �����  �           ����    6 7          � � �� r     5  Lm  ܌   ��  �       ��b       ���� � �����  �           ����    8 9          � �� s     d  �n  $�   ��  �       ��b       ���� � �����  �           ����    ; <          � 	�� t     �  p  l�   ��  �       ��b       ����  �����  �           ����    = >          � �� u     �  �q  ��   ��  �       ��b       ���� �����  �           ����    ? @          � �� v     �  �r  ��   ��  �       ��b       ���� �����  �           ����    A B          � �� w       Tt  D�   ��  �	       ��b       ���� A  �  �           ����    2 3          � �� x       �y  X�      �        ��c        ���� � �����  �           ����    4 5          � 	�� y     I  z{  ��       �       ��c        ���� � �����  �           ����    6 7          � �� z     �   }   �   ��  �       ��c        ���� � �����  �           ����    8 9          � �� {     �  �~  T�   ��  �       ��c       ���� � �����  �           ����    : ;          � �� |     �  �  �    ��  �       ��c       ����  �����  �           ����    < =          � !�� }     #  ��  �   ��  �       ��c       ���� �����  �           ����    ? @          � '�� ~     Z  �  P+   ��  �       ��c       ���� �����  �           ����    A B          � -�      �  ��  �@   ��  �       ��c       ���� �����  �           ����    C D          � 3	� �     �  $�  �U   ��  �       ��c       ���� �����  �           ����    E F          � 9� �     �  ��  Lk   ��  �	       ��c       ���� #K  �  �            ����                             ,  h       �        ��d        ���� � ������������          ����                 "            J  �       �       ��d        ���� � ������������          ����                 '            h  �       �       ��d        ���� � ������������          ����                 ,            �         �       ��d       ���� � ������������          ����   	 
             1            �  H       �       ��d       ���� � ������������          ����                 6         	   �  �       �       ��d       ���� � ������������          ����                 ;         	   �  �       �       ��d       ���� � ������������          ����                 @         
   �  �       �       ��d       ���� � ������������          ����                 E         
     8       �       ��d       ���� � ������������          ����                 J            :  t       �	       ��d       ���� � ������������          ����                $ 8            �         �        ��e        ���� � ������������          ����                ' =            �  �       �       ��e        ���� � ������������          ����   	 
            * B            *  ~	       �       ��e        ���� � ������������          ����                - G            f  2
       �       ��e       ���� � ������������          ����                0 L            �  �
       �       ��e       ���� � ������������          ����                3 Q            �  �       �       ��e       ���� � ������������          ����                6 V              N       �       ��e       ���� � ������������          ����                9 [         !   V         �       ��e       ���� � ������������          ����                < `         #   �  �       �       ��e       ���� � ������������          ����                ? e         $   �  j       �	       ��e       ���� � ������������          ����   	 
           + R         :   �  �       �        ��f        ���� � ������������         ����              ! / W         >     `       �       ��f        ���� � ������������         ����              $ 3 \         B   r  �       �       ��f        ���� � ������������         ����              ' 7 a         E   �  0       �       ��f       ���� � ������������         ����              * ; f         I   &  �       �       ��f       ���� � ������������         ����              - ? k         L   �          �       ��f       ���� � ������������         ����              0 C p         P   �  h       �       ��f       ���� � ������������         ����              3 G u         T   4  �        �       ��f       ���� � ������������         ����              6 K z         W   �  8"       �       ��f       ���� � ������������         ����              9 O          [   �  �#       �	       ��f       ���� � ������������          ����              & < k        �   P
  �3       �        ��g        ���� � ������������         ����              ) @ q        �   �
  �5       �       ��g        ���� � ������������         ����              , D w         �   @  @8       �       ��g        ���� � ������������         ����              / H } #       �   �  �:       �       ��g       ���� � ������������         ����              2 L � &       �   0  �<       �       ��g       ���� � ������������         ����              5 P � )       �   �  H?       �       ��g       ���� � ������������         ����              8 T � ,       �      �A       �       ��g       ���� � ������������         ����              ; X � /       �   �  �C       �       ��g       ���� � ������������         ����              > \ � 2       �     PF       �       ��g       ���� � ������������         ����     !          A ` � 5       �   �  �H       �	       ��g       ���� � ������������          ����              - L � !       �   h  pb       �        ��h        ���� � ������������         ����              0 P � $         �  �e       �       ��h        ���� � ������������         ����              3 T � '         �  xi       �       ��h        ���� � ������������         ����              6 X � *         *  �l       �       ��h       ���� � ������������         ����              9 \ � -          �  �p       �       ��h       ���� � ������������         ����              < ` � 0       )  V  t       �       ��h       ���� � ������������         ����              ? d � 3       2  �  �w       �       ��h       ���� � ������������         ����     !          B h � 6       ;  �  {       �       ��h       ���� � ������������         ����   " #          E l � 9       D    �~    
   �       ��h       ���� � ������������         ����   $ %          H p � <       M  �  �    	   �	       ��h       ���� � ������������          ����              4 [ � (       �    *�       �        ��i        ���� � ������������         ����              8 _ � +       �  �  �       �       ��i        ���� � ������������         ����              < c � .       �  n  �       �       ��i        ���� � ������������         ����              @ g � 1       �  "  �       �       ��i       ���� � ������������         ����              D k � 4       �  �  ڻ       �       ��i       ���� � ������������         ����     !          H o � 7       �  �  ��       �       ��i       ���� � ������������         ����   " #          L s � :       �  >  ��       �       ��i       ���� � ������������         ����   $ %          P w � =         �  ��    	   �       ��i       ���� � ������������         ����   & '          T { � @         �  ��       �       ��i       ���� � ������������         ����   ( )          X  � C         Z  v�       �	       ��i       ���� � ������������         ����              D j � .       �  *!  P	      �        ��j        ���� � �����  �           ����              H o � 2       �  �!  �      �       ��j        ���� � �����  �           ����              L t � 6       �  �"  p      �       ��j        ���� � �����  �           ����               P y � :       �  �#         �       ��j       ���� � �����  �           ����   ! "          T ~ � >       �  r$  �#      �       ��j       ���� � �����  �           ����   $ %          X � � B       �  D%   *   	   �       ��j       ���� � �����  �           ����   & '          \ � � F         &  �0      �       ��j       ���� � �����  �           ����   ( )          ` � � J         �&  @7      �       ��j       ���� � �����  �           ����   * +          d �  N       -  �'  �=      �       ��j       ���� � �����  �           ����   , -          h � R       >  �(  `D      �	       ��j       ���� � �����  �           ����              T � � >       �  �+  t�      �        ��k        ���� � �����  �           ����               X � � B         �,  �      �       ��k        ���� � �����  �           ����   ! "          \ � � F         �-  T�      �       ��k        ���� � �����  �           ����   # $          ` � J       2  �.  ģ   	   �       ��k       ���� � �����  �           ����   % &          d � N       H  �/  4�      �       ��k       ���� � �����  �           ����   ' (          h � R       ]  �0  ��      �       ��k       ���� � �����  �           ����   * +          l � V       s  t1  �      �       ��k       ���� � �����  �           ����   , -          p � !Z       �  d2  ��      �       ��k       ���� � �����  �           ����   . /          t � (^       �  T3  ��      �       ��k       ���� � �����  �           ����   0 1          x � /b       �  D4  d�      �	       ��k       ���� � -  �  �           ����   ! "          c � M       �  8  (0      �      	  ��l        ����	 � �����  �           ����   # $          g �  Q       �  9  �:   
   �     	  ��l        ����	 � �����  �           ����   % &          k � 'U       �   :  @E      �     	  ��l        ����	 � �����  �           ����   ' (          o � .Y       �  .;  �O      �     	  ��l       ����	 � �����  �           ����   ) *          s � 5]         <<  XZ      �     	  ��l       ����	 � �����  �           ����   + ,          w � <a       !  J=  �d      �     	  ��l       ����	 � �����  �           ����   . /          { � Ce       <  X>  po      �     	  ��l       ����	 � �����  �           ����   0 1           � Ji       W  f?  �y      �     	  ��l       ����	 � �����  �           ����   2 3          � � Qm       r  t@  ��       �     	  ��l       ����	 � �����  �           ����   4 5          � � Xq       �  �A  �   ��  �	     	  ��l       ����	 � 7  �  �           ����   % &          r � A\       �  �E  ��   	   �      
  ��m        ����
 � �����  �           ����   ' (          w � H`       �  �F  �      �     
  ��m        ����
 � �����  �           ����   ) *          | � Od       �  H  �      �     
  ��m        ����
 � �����  �           ����   + ,          � � Vh         >I  �%      �     
  ��m       ����
 � �����  �           ����   - .          � � ]l       /  jJ  �2      �     
  ��m       ����
 � �����  �           ����   / 0          � � dp       P  �K  r?      �     
  ��m       ����
 � �����  �           ����   2 3          � � kt       q  �L  VL      �     
  ��m       ����
 � �����  �           ����   4 5          � � rx       �  �M  :Y   ��  �     
  ��m       ����
 � �����  �           ����   6 7          � � y|       �  O  f   ��  �     
  ��m       ����
 � �����  �           ����   8 9          � � ��       �  FP  s   ��  �	     
  ��m       ����
 7  �  �           ����   ) *          � � hj d     2
  �T  ��      �        ��n        ���� � �����  �           ����   + ,          � � oo e     Y
  @V         �       ��n        ���� � �����  �           ����   - .          � � vt f     �
  �W  x      �       ��n        ���� � �����  �           ����   / 0          � � }y g     �
  �X  �)      �       ��n       ���� � �����  �           ����   1 2          � � �~ h     �
  Z  h9      �       ��n       ���� � �����  �           ����   3 4          � � �� i     �
  h[  �H   ��  �       ��n       ���� � �����  �           ����   6 7          � � �� j       �\  XX   ��  �       ��n       ���� � �����  �           ����   8 9          � � �� k     G  �]  �g   ��  �       ��n       ���� � �����  �           ����   : ;          � � �� l     n  F_  Hw   ��  �       ��n       ���� �����  �           ����   < =          � � �� m     �  �`  ��   ��  �	       ��n       ���� A  �  �           ����   - .          � � �� n     9  �e  X*      �        ��o        ���� � �����  �           ����   / 0          � � �� o     h   g  �<      �       ��o        ���� � �����  �           ����   1 2          � � �� p     �  �h  �N      �       ��o        ���� � �����  �           ����   3 4          � � �� q     �  �i  0a   ��  �       ��o       ���� � �����  �           ����   5 6          � � �� r     �  Xk  xs   ��  �       ��o       ���� � �����  �           ����   7 8          � �� s     #  �l  ��   ��  �       ��o       ���� � �����  �           ����   : ;          � 	�� t     R  (n  �   ��  �       ��o       ����  �����  �           ����   < =          � �� u     �  �o  P�   ��  �       ��o       ���� �����  �           ����   > ?          � �� v     �  �p  ��   ��  �       ��o       ���� �����  �           ����   @ A          � �� w     �  `r  ��   ��  �	       ��o       ���� A  �  �           ����   1 2          � �� x     �   x   �      �        ��p        ���� � �����  �           ����   3 4          � 	�� y       �y  T�       �       ��p        ���� � �����  �           ����   5 6          � �� z     :  {  ��   ��  �       ��p        ���� � �����  �           ����   7 8          � �� {     p  �|  ��   ��  �       ��p       ���� � �����  �           ����   9 :          � �� |     �  ~  P�   ��  �       ��p       ����  �����  �           ����   ; <          � !�� }     �  �  ��   ��  �       ��p       ���� �����  �           ����   > ?          � '�� ~       $�  �   ��  �       ��p       ���� �����  �           ����   @ A          � -��      K  ��  L%   ��  �       ��p       ���� �����  �           ����   B C          � 3�� �     �  0�  �:   ��  �       ��p       ���� �����  �           ����   D E          � 9� �     �  ��  �O   ��  �	       ��p       ���� #K  �  �            ����                % %            �   �        E        ��q        ���� � ������������          ����                % *            �   �       E       ��q        ���� � ������������          ����                % /                     E       ��q        ���� � ������������          ����                % 4            "  D       E       ��q       ���� � ������������          ����   	 
            % 9            @  �       E       ��q       ���� � ������������          ����                % >            ^  �       E       ��q       ���� � ������������          ����                % C            |  �       E       ��q       ���� � ������������          ����                % H            �  4       E       ��q       ���� � ������������          ����                % M            �  p       E       ��q       ���� � ������������          ����                % R         	   �  �       E	       ��q       ���� � ������������          ����                $ @            N  �       F        ��r        ���� � ������������          ����                ' E            �  �       F       ��r        ���� � ������������          ����   	 
            * J            �  R       F       ��r        ���� � ������������          ����                - O              	       F       ��r       ���� � ������������          ����                0 T            >  �	       F       ��r       ���� � ������������          ����                3 Y            z  n
       F       ��r       ���� � ������������          ����                6 ^            �  "       F       ��r       ���� � ������������          ����                9 c            �  �       F       ��r       ���� � ������������          ����                < h             .  �       F       ��r       ���� � ������������          ����                ? m         !   j  >       F	       ��r       ���� � ������������         ����   	 
           + Z         6   Z  h       G        ��s        ���� � ������������         ����              ! / _         :   �  �       G       ��s        ���� � ������������         ����              $ 3 d         >     8       G       ��s        ���� � ������������         ����              ' 7 i         A   h  �       G       ��s       ���� � ������������         ����              * ; n         E   �         G       ��s       ���� � ������������         ����              - ? s         H     p       G       ��s       ���� � ������������         ����              0 C x         L   v  �       G       ��s       ���� � ������������         ����              3 G }         P   �  @       G       ��s       ���� � ������������         ����              6 K �         S   *  �        G       ��s       ���� � ������������         ����              9 O �         W   �  "       G	       ��s       ���� � ������������         ����              & < s           �	  �1       H        ��t        ���� � ������������          ����              ) @ y        �   d
  �3       H       ��t        ���� � ������������          ����              , D          �   �
  L6       H       ��t        ���� � ������������          ����              / H � #       �   T  �8       H       ��t       ���� � ������������          ����              2 L � &       �   �  �:       H       ��t       ���� � ������������          ����              5 P � )       �   D  T=       H       ��t       ���� � ������������          ����              8 T � ,       �   �  �?       H       ��t       ���� � ������������          ����              ; X � /       �   4  B       H       ��t       ���� � ������������          ����              > \ � 2       �   �  \D       H       ��t       ���� � ������������          ����     !          A ` � 5       �   $  �F       H	       ��t       ���� � ������������          ����              - L � !       �     `       I        ��u        ���� � ������������!         ����              0 P � $       �   �  �c       I       ��u        ���� � ������������!         ����              3 T � '         0   g       I       ��u        ���� � ������������!         ����              6 X � *         �  �j       I       ��u       ���� � ������������!         ����              9 \ � -         \  (n       I       ��u       ���� � ������������!         ����              < ` � 0       #  �  �q       I       ��u       ���� � ������������!         ����              ? d � 3       ,  �  0u       I       ��u       ���� � ������������!         ����     !          B h � 6       5    �x       I       ��u       ���� � ������������!         ����   " #          E l � 9       >  �  8|    
   I       ��u       ���� � ������������!         ����   $ %          H p � <       G  J  �    	   I	       ��u       ���� � ������������!         ����              4 [ � (       �  �  n�       J        ��v        ���� � ������������"         ����              8 _ � +       �  V  Z�       J       ��v        ���� � ������������"         ����              < c � .       �  
  F�       J       ��v        ���� � ������������"         ����              @ g � 1       �  �  2�       J       ��v       ���� � ������������"         ����              D k � 4       �  r  �       J       ��v       ���� � ������������"         ����     !          H o � 7       �  &  
�       J       ��v       ���� � ������������"         ����   " #          L s � :       �  �  ��       J       ��v       ���� � ������������"         ����   $ %          P w � =       �  �  ��    	   J       ��v       ���� � ������������"         ����   & '          T { � @         B  ��       J       ��v       ���� � ������������"         ����   ( )          X  � C         �  ��       J	       ��v       ���� � ������������"         ����              D j � .       �  �   0      K        ��w        ���� � �����  �  #         ����              H o � 2       �  �!  �      K       ��w        ���� � �����  �  #         ����              L t � 6       �  j"  P      K       ��w        ���� � �����  �  #         ����               P y � :       �  <#  �      K       ��w       ���� � �����  �  #         ����   ! "          T ~ � >       �  $  p       K       ��w       ���� � �����  �  #         ����   $ %          X � � B       �  �$   '   	   K       ��w       ���� � �����  �  #         ����   & '          \ � � F         �%  �-      K       ��w       ���� � �����  �  #         ����   ( )          ` � J         �&   4      K       ��w       ���� � �����  �  #         ����   * +          d � N       %  V'  �:      K       ��w       ���� � �����  �  #         ����   , -          h � R       6  ((  @A      K	       ��w       ���� � �����  �  #         ����              T � � >       �  p+  ��      L        ��x        ���� � �����  �  $         ����               X � � B       �  `,  `�      L       ��x        ���� � �����  �  $         ����   ! "          \ � F         P-  З      L       ��x        ���� � �����  �  $         ����   # $          ` � J       )  @.  @�   	   L       ��x       ���� � �����  �  $         ����   % &          d � N       ?  0/  ��      L       ��x       ���� � �����  �  $         ����   ' (          h � R       T   0   �      L       ��x       ���� � �����  �  $         ����   * +          l � "V       j  1  ��      L       ��x       ���� � �����  �  $         ����   , -          p � )Z       �   2   �      L       ��x       ���� � �����  �  $         ����   . /          t � 0^       �  �2  p�      L       ��x       ���� � �����  �  $         ����   0 1          x � 7b       �  �3  ��      L	       ��x       ���� � -  �  �  $         ����   ! "          c � !M       �  �7  @,      M      	  ��y        ����	 � �����  �  %         ����   # $          g � (Q       �  �8  �6   
   M     	  ��y        ����	 � �����  �  %         ����   % &          k � /U       �  �9  XA      M     	  ��y        ����	 � �����  �  %         ����   ' (          o � 6Y       �  �:  �K      M     	  ��y       ����	 � �����  �  %         ����   ) *          s � =]       �  �;  pV      M     	  ��y       ����	 � �����  �  %         ����   + ,          w � Da         �<  �`      M     	  ��y       ����	 � �����  �  %         ����   . /          { � Ke       2  �=  �k      M     	  ��y       ����	 � �����  �  %         ����   0 1           � Ri       M  ?  v      M     	  ��y       ����	 � �����  �  %         ����   2 3          � � Ym       h  @  ��       M     	  ��y       ����	 � �����  �  %         ����   4 5          � � `q       �  A  ,�   ��  M	     	  ��y       ����	 � 7  �  �  %         ����   % &          r � I\       �  VE  ��   	   N      
  ��z        ����
 � �����  �  &         ����   ' (          w � P`       �  �F  �      N     
  ��z        ����
 � �����  �  &         ����   ) *          | � Wd       �  �G  z      N     
  ��z        ����
 � �����  �  &         ����   + ,          � � ^h         �H  ^!      N     
  ��z       ����
 � �����  �  &         ����   - .          � � el       $  J  B.      N     
  ��z       ����
 � �����  �  &         ����   / 0          � � lp       E  2K  &;      N     
  ��z       ����
 � �����  �  &         ����   2 3          � � st       f  ^L  
H      N     
  ��z       ����
 � �����  �  &         ����   4 5          � � zx       �  �M  �T   ��  N     
  ��z       ����
 � �����  �  &         ����   6 7          � � �|       �  �N  �a   ��  N     
  ��z       ����
 � �����  �  &         ����   8 9          � � ��       �  �O  �n   ��  N	     
  ��z       ����
 7  �  �  &         ����   ) *          � � pj d     &
  �T  ��      O        ��{        ���� � �����  �  '         ����   + ,          � � wo e     M
  �U  P      O       ��{        ���� � �����  �  '         ����   - .          � � ~t f     u
  &W  �      O       ��{        ���� � �����  �  '         ����   / 0          � � �y g     �
  pX  @%      O       ��{       ���� � �����  �  '         ����   1 2          � � �~ h     �
  �Y  �4      O       ��{       ���� � �����  �  '         ����   3 4          � � �� i     �
  [  0D   ��  O       ��{       ���� � �����  �  '         ����   6 7          � � �� j       N\  �S   ��  O       ��{       ���� � �����  �  '         ����   8 9          � � �� k     ;  �]   c   ��  O       ��{       ���� � �����  �  '         ����   : ;          � � �� l     b  �^  �r   ��  O       ��{       ���� �����  �  '         ����   < =          � � �� m     �  ,`  �   ��  O	       ��{       ���� A  �  �  '         ����   - .          � � �� n     ,  Te  D%      P        ��|        ���� � �����  �  (         ����   / 0          � � �� o     [  �f  �7      P       ��|        ���� � �����  �  (         ����   1 2          � � �� p     �  $h  �I      P       ��|        ���� � �����  �  (         ����   3 4          � � �� q     �  �i  \   ��  P       ��|       ���� � �����  �  (         ����   5 6          � � �� r     �  �j  dn   ��  P       ��|       ���� � �����  �  (         ����   7 8          � �� s       \l  ��   ��  P       ��|       ���� � �����  �  (         ����   : ;          � 	�� t     E  �m  ��   ��  P       ��|       ����  �����  �  (         ����   < =          � �� u     s  ,o  <�   ��  P       ��|       ���� �����  �  (         ����   > ?          � �� v     �  �p  ��   ��  P       ��|       ���� �����  �  (         ����   @ A          � �� w     �  �q  ��   ��  P	       ��|       ���� A  �  �  (         ����   1 2          � �� x     �  �w  ��      Q        ��}        ���� � �����  �  )         ����   3 4          � 	�� y     �  "y  ܟ       Q       ��}        ���� � �����  �  )         ����   5 6          � �� z     ,  �z  0�   ��  Q       ��}        ���� � �����  �  )         ����   7 8          � �� {     b  .|  ��   ��  Q       ��}       ���� � �����  �  )         ����   9 :          � �� |     �  �}  ��   ��  Q       ��}       ����  �����  �  )         ����   ; <          � !�� }     �  :  ,�   ��  Q       ��}       ���� �����  �  )         ����   > ?          � '�� ~       ��  �
   ��  Q       ��}       ���� �����  �  )         ����   @ A          � -��      =  F�  �   ��  Q       ��}       ���� �����  �  )         ����   B C          � 3� �     s  ̃  (5   ��  Q       ��}       ���� �����  �  )         ����   D E          � 9� �     �  R�  |J   ��  Q	       ��}       ���� #K  �  �  )          ����                          !   �  /       �        ��~        ���� � ������������*          ����                          (   �  �       �       ��~        ���� � ������������*          ����                 #         )            �       ��~        ���� � ������������*          ����                 (         )   *  T       �       ��~       ���� � ������������*          ����   	 
             -         *   H  �       �       ��~       ���� � ������������*          ����                 2         +   f  �       �       ��~       ���� � ������������*          ����                 7         +   �         �       ��~       ���� � ������������*          ����                 <         ,   �  D       �       ��~       ���� � ������������*          ����                 A         ,   �  �       �       ��~       ���� � ������������*          ����                 F         -   �  �       �	       ��~       ���� � ������������*          ����                $ 4         G   V	         �        ��        ���� � ������������+          ����                ' 9         I   �	  �       �       ��        ���� � ������������+          ����   	 
            * >         K   �	  j       �       ��        ���� � ������������+          ����                - C         M   

         �       ��       ���� � ������������+          ����                0 H         N   F
  �       �       ��       ���� � ������������+          ����                3 M         P   �
  �       �       ��       ���� � ������������+          ����                6 R         R   �
  :        �       ��       ���� � ������������+          ����                9 W         T   �
  �        �       ��       ���� � ������������+          ����                < \         V   6  �!       �       ��       ���� � ������������+          ����                ? a         W   r  V"       �	       ��       ���� � ������������+          ����   	 
           + N         ~   b  �1       �        ���        ���� � ������������,         ����              ! / S         �   �  �2       �       ���        ���� � ������������,         ����              $ 3 X         �     X4       �       ���        ���� � ������������,         ����              ' 7 ]         �   p  �5       �       ���       ���� � ������������,         ����              * ; b         �   �  (7       �       ���       ���� � ������������,         ����              - ? g         �   $  �8       �       ���       ���� � ������������,         ����              0 C l         �   ~  �9       �       ���       ���� � ������������,         ����              3 G q         �   �  `;       �       ���       ���� � ������������,         ����              6 K v         �   2  �<       �       ���       ���� � ������������,         ����              9 O {         �   �  0>       �	       ���       ���� � ������������,          ����              & < g        �   �  �T       �        ���        ���� � ������������-         ����              ) @ m        �   l  W       �       ���        ���� � ������������-         ����              , D s         �   �  tY       �       ���        ���� � ������������-         ����              / H y #       �   \  �[       �       ���       ���� � ������������-         ����              2 L  &       �   �  $^       �       ���       ���� � ������������-         ����              5 P � )       �   L  |`       �       ���       ���� � ������������-         ����              8 T � ,       �   �  �b       �       ���       ���� � ������������-         ����              ; X � /         <  ,e       �       ���       ���� � ������������-         ����              > \ � 2       	  �  �g       �       ���       ���� � ������������-         ����     !          A ` � 5         ,  �i       �	       ���       ���� � ������������-          ����              - L � !       b    H�       �        ���        ���� � ������������.         ����              0 P � $       k  �  ̍       �       ���        ���� � ������������.         ����              3 T � '       t  8  P�       �       ���        ���� � ������������.         ����              6 X � *       }  �  Ԕ       �       ���       ���� � ������������.         ����              9 \ � -       �  d  X�       �       ���       ���� � ������������.         ����              < ` � 0       �  �  ܛ       �       ���       ���� � ������������.         ����              ? d � 3       �  �  `�       �       ���       ���� � ������������.         ����     !          B h � 6       �  &  �       �       ���       ���� � ������������.         ����   " #          E l � 9       �  �  h�    
   �       ���       ���� � ������������.         ����   $ %          H p � <       �  R  �    	   �	       ���       ���� � ������������.          ����              4 [ � (       %  �  ��       �        ���        ���� � ������������/         ����              8 _ � +       2  ^  ��       �       ���        ���� � ������������/         ����              < c � .       >     ~�       �       ���        ���� � ������������/         ����              @ g � 1       K  �   j�       �       ���       ���� � ������������/         ����              D k � 4       W  z!  V�       �       ���       ���� � ������������/         ����     !          H o � 7       d  ."  B�       �       ���       ���� � ������������/         ����   " #          L s � :       q  �"  .�       �       ���       ���� � ������������/         ����   $ %          P w � =       }  �#  �    	   �       ���       ���� � ������������/         ����   & '          T { � @       �  J$  �       �       ���       ���� � ������������/         ����   ( )          X  � C       �  �$  �      �	       ���       ���� � ������������/         ����              D j � .       /  �'  p>      �        ���        ���� � �����  �  0         ����              H o � 2       @  �(   E      �       ���        ���� � �����  �  0         ����              L t � 6       P  r)  �K      �       ���        ���� � �����  �  0         ����               P y � :       a  D*   R      �       ���       ���� � �����  �  0         ����   ! "          T ~ � >       r  +  �X      �       ���       ���� � �����  �  0         ����   $ %          X � � B       �  �+  @_   	   �       ���       ���� � �����  �  0         ����   & '          \ � � F       �  �,  �e      �       ���       ���� � �����  �  0         ����   ( )          ` � � J       �  �-  `l      �       ���       ���� � �����  �  0         ����   * +          d � � N       �  ^.  �r      �       ���       ���� � �����  �  0         ����   , -          h � R       �  0/  �y      �	       ���       ���� � �����  �  0         ����              T � � >       �  x2  8�      �        ���        ���� � �����  �  1         ����               X � � B       �  h3  ��      �       ���        ���� � �����  �  1         ����   ! "          \ � � F       �  X4  �      �       ���        ���� � �����  �  1         ����   # $          ` � J       �  H5  ��   	   �       ���       ���� � �����  �  1         ����   % &          d � N       �  86  ��      �       ���       ���� � �����  �  1         ����   ' (          h � R       �  (7  h�      �       ���       ���� � �����  �  1         ����   * +          l � V         8  ��      �       ���       ���� � �����  �  1         ����   , -          p � Z       "  9  H      �       ���       ���� � �����  �  1         ����   . /          t � $^       7  �9  �	      �       ���       ���� � �����  �  1         ����   0 1          x � +b       M  �:  (      �	       ���       ���� � -  �  �  1         ����   ! "          c � M       D  �>  �r      �      	  ���        ����	 � �����  �  2         ����   # $          g � Q       _  �?  }   
   �     	  ���        ����	 � �����  �  2         ����   % &          k � #U       z  �@  ��      �     	  ���        ����	 � �����  �  2         ����   ' (          o � *Y       �  �A  4�      �     	  ���       ����	 � �����  �  2         ����   ) *          s � 1]       �  �B  ��      �     	  ���       ����	 � �����  �  2         ����   + ,          w � 8a       �  �C  L�      �     	  ���       ����	 � �����  �  2         ����   . /          { � ?e       �  �D  ر      �     	  ���       ����	 � �����  �  2         ����   0 1           � Fi         
F  d�      �     	  ���       ����	 � �����  �  2         ����   2 3          � � Mm         G  ��       �     	  ���       ����	 � �����  �  2         ����   4 5          � � Tq       7  &H  |�   ��  �	     	  ���       ����	 � 7  �  �  2         ����   % &          r � =\       f  ^L  
H   	   �      
  ���        ����
 � �����  �  3         ����   ' (          w � D`       �  �M  �T      �     
  ���        ����
 � �����  �  3         ����   ) *          | � Kd       �  �N  �a      �     
  ���        ����
 � �����  �  3         ����   + ,          � � Rh       �  �O  �n      �     
  ���       ����
 � �����  �  3         ����   - .          � � Yl       �  Q  �{      �     
  ���       ����
 � �����  �  3         ����   / 0          � � `p       	  :R  ~�      �     
  ���       ����
 � �����  �  3         ����   2 3          � � gt       ,	  fS  b�      �     
  ���       ����
 � �����  �  3         ����   4 5          � � nx       M	  �T  F�   ��  �     
  ���       ����
 � �����  �  3         ����   6 7          � � u|       n	  �U  *�   ��  �     
  ���       ����
 � �����  �  3         ����   8 9          � � |�       �	  �V  �   ��  �	     
  ���       ����
 7  �  �  3         ����   ) *          � � dj d     �
  �[  8K      �        ���        ���� � �����  �  4         ����   + ,          � � ko e     %  �\  �Z      �       ���        ���� � �����  �  4         ����   - .          � � rt f     M  .^  (j      �       ���        ���� � �����  �  4         ����   / 0          � � yy g     t  x_  �y      �       ���       ���� � �����  �  4         ����   1 2          � � �~ h     �  �`  �      �       ���       ���� � �����  �  4         ����   3 4          � � �� i     �  b  ��   ��  �       ���       ���� � �����  �  4         ����   6 7          � � �� j     �  Vc  �   ��  �       ���       ���� � �����  �  4         ����   8 9          � � �� k       �d  ��   ��  �       ���       ���� � �����  �  4         ����   : ;          � � �� l     :  �e  ��   ��  �       ���       ���� �����  �  4         ����   < =          � � �� m     b  4g  p�   ��  �	       ���       ���� A  �  �  4         ����   - .          � � �� n       \l  ��      �        ���        ���� � �����  �  5         ����   / 0          � � �� o     E  �m  ��      �       ���        ���� � �����  �  5         ����   1 2          � � �� p     s  ,o  <�      �       ���        ���� � �����  �  5         ����   3 4          � � �� q     �  �p  ��   ��  �       ���       ���� � �����  �  5         ����   5 6          � � �� r     �  �q  ��   ��  �       ���       ���� � �����  �  5         ����   7 8          � �� s        ds  �   ��  �       ���       ���� � �����  �  5         ����   : ;          � 	�� t     /  �t  \�   ��  �       ���       ����  �����  �  5         ����   < =          � �� u     ]  4v  �    ��  �       ���       ���� �����  �  5         ����   > ?          � �� v     �  �w  �   ��  �       ���       ���� �����  �  5         ����   @ A          � �� w     �  y  4%   ��  �	       ���       ���� A  �  �  5         ����   1 2          � �� x     �  �~  ��      �        ���        ���� � �����  �  6         ����   3 4          � 	�� y     �  *�  L       �       ���        ���� � �����  �  6         ����   5 6          � �� z     (  ��  �   ��  �       ���        ���� � �����  �  6         ����   7 8          � �� {     ^  6�  �,   ��  �       ���       ���� � �����  �  6         ����   9 :          � �� |     �  ��  HB   ��  �       ���       ����  �����  �  6         ����   ; <          � !�� }     �  B�  �W   ��  �       ���       ���� �����  �  6         ����   > ?          � '�� ~       ȇ  �l   ��  �       ���       ���� �����  �  6         ����   @ A          � -��      9  N�  D�   ��  �       ���       ���� �����  �  6         ����   B C          � 3�� �     o  Ԋ  ��   ��  �       ���       ���� �����  �  6         ����   D E          � 9� �     �  Z�  �   ��  �	       ���       ���� #K  �  �  6          ����                1 1            @  �                ���        ���� � ������������7          ����                1 6             ^  �               ���        ���� � ������������7          ����                1 ;         !   |  �               ���        ���� � ������������7          ����    	            1 @         !   �  4               ���       ���� � ������������7          ����   
             1 E         "   �  p               ���       ���� � ������������7          ����                1 J         #   �  �               ���       ���� � ������������7          ����                1 O         #   �  �               ���       ���� � ������������7          ����                1 T         $     $               ���       ���� � ������������7          ����                1 Y         $   0  `               ���       ���� � ������������7          ����                1 ^         %   N  �       	        ���       ���� � ������������7          ����                $ L         ;   �  R               ���        ���� � ������������8          ����    	            ' Q         =                   ���        ���� � ������������8          ����   
             * V         ?   >  �              ���        ���� � ������������8          ����                - [         A   z  n              ���       ���� � ������������8          ����                0 `         B   �  "              ���       ���� � ������������8          ����                3 e         D   �  �              ���       ���� � ������������8          ����                6 j         F   .	  �              ���       ���� � ������������8          ����                9 o         H   j	  >              ���       ���� � ������������8          ����                < t         J   �	  �              ���       ���� � ������������8          ����                ? y         K   �	  �       	       ���       ���� � ������������8         ����   
            + f         n   �
  H+               ���        ���� � ������������9         ����              ! / k         r   ,  �,              ���        ���� � ������������9         ����              $ 3 p         v   �  .              ���        ���� � ������������9         ����              ' 7 u         y   �  �/              ���       ���� � ������������9         ����              * ; z         }   :  �0              ���       ���� � ������������9         ����              - ?          �   �  P2              ���       ���� � ������������9         ����              0 C �         �   �  �3              ���       ���� � ������������9         ����              3 G �         �   H   5              ���       ���� � ������������9         ����              6 K �         �   �  �6              ���       ���� � ������������9         ����              9 O �         �   �  �7       	       ���       ���� � ������������9         ����              & <         �   d  �L               ���        ���� � ������������:         ����              ) @ �        �   �  LO              ���        ���� � ������������:         ����              , D �         �   T  �Q              ���        ���� � ������������:         ����              / H � #       �   �  �S              ���       ���� � ������������:         ����              2 L � &       �   D  TV              ���       ���� � ������������:         ����              5 P � )       �   �  �X              ���       ���� � ������������:         ����              8 T � ,       �   4  [              ���       ���� � ������������:         ����              ; X � /       �   �  \]              ���       ���� � ������������:         ����               > \ � 2       �   $  �_              ���       ���� � ������������:         ����   ! "          A ` � 5       �   �  b       	       ���       ���� � ������������:         ����              - L � !       J  |  �               ���        ���� � ������������;         ����              0 P � $       S    l�              ���        ���� � ������������;         ����              3 T � '       \  �  ��              ���        ���� � ������������;         ����              6 X � *       e  >  t�              ���       ���� � ������������;         ����              9 \ � -       n  �  ��              ���       ���� � ������������;         ����              < ` � 0       w  j  |�              ���       ���� � ������������;         ����               ? d � 3       �      �              ���       ���� � ������������;         ����   ! "          B h � 6       �  �  ��              ���       ���� � ������������;         ����   # $          E l � 9       �  ,  �    
          ���       ���� � ������������;         ����   % &          H p � <       �  �  ��    	   	       ���       ���� � ������������;         ����              4 [ � (       	    ��               ���        ���� � ������������<         ����              8 _ � +         �  ��              ���        ���� � ������������<         ����              < c � .       "  �  ��              ���        ���� � ������������<         ����              @ g � 1       /  6  z�              ���       ���� � ������������<         ����              D k � 4       ;  �  f�              ���       ���� � ������������<         ����   ! "          H o � 7       H  �   R�              ���       ���� � ������������<         ����   # $          L s � :       U  R!  >�              ���       ���� � ������������<         ����   % &          P w � =       a  "  *�    	          ���       ���� � ������������<         ����   ' (          T { � @       n  �"  �              ���       ���� � ������������<         ����   ) *          X  � C       z  n#  �       	       ���       ���� � ������������<         ����              D j � .         >&  �1              ���        ���� � �����  �  =         ����              H o � 2          '  �8             ���        ���� � �����  �  =         ����              L t � 6       0  �'  ?             ���        ���� � �����  �  =         ����     !          P y � :       A  �(  �E             ���       ���� � �����  �  =         ����   " #          T ~ � >       R  �)  0L             ���       ���� � �����  �  =         ����   $ %          X � B       c  X*  �R   	          ���       ���� � �����  �  =         ����   ' (          \ � F       t  *+  PY             ���       ���� � �����  �  =         ����   ) *          ` � J       �  �+  �_             ���       ���� � �����  �  =         ����   + ,          d � N       �  �,  pf             ���       ���� � �����  �  =         ����   - .          h � R       �  �-   m      	       ���       ���� � �����  �  =         ����              T � >       f  �0  (�              ���        ���� � �����  �  >         ����     !          X � B       |  �1  ��             ���        ���� � �����  �  >         ����   " #          \ � F       �  �2  �             ���        ���� � �����  �  >         ����   $ %          ` � J       �  �3  x�   	          ���       ���� � �����  �  >         ����   & '          d �  N       �  �4  ��             ���       ���� � �����  �  >         ����   ( )          h � 'R       �  �5  X�             ���       ���� � �����  �  >         ����   + ,          l � .V       �  �6  ��             ���       ���� � �����  �  >         ����   - .          p � 5Z       �  x7  8�             ���       ���� � �����  �  >         ����   / 0          t � <^         h8  ��             ���       ���� � �����  �  >         ����   1 2          x � Cb       )  X9        	       ���       ���� � -  �  �  >         ����   " #          c � -M         =  �b              ���        ����	 � �����  �  ?         ����   $ %          g � 4Q       7  &>  |m   
          ���        ����	 � �����  �  ?         ����   & '          k � ;U       R  4?  x             ���        ����	 � �����  �  ?         ����   ( )          o � BY       m  B@  ��             ���       ����	 � �����  �  ?         ����   * +          s � I]       �  PA   �             ���       ����	 � �����  �  ?         ����   , -          w � Pa       �  ^B  ��             ���       ����	 � �����  �  ?         ����   / 0          { � We       �  lC  8�             ���       ����	 � �����  �  ?         ����   1 2           � ^i       �  zD  Ĭ             ���       ����	 � �����  �  ?         ����   3 4          � � em       �  �E  P�              ���       ����	 � �����  �  ?         ����   5 6          � � lq         �F  ��   ��  	       ���       ����	 � 7  �  �  ?         ����   & '          r � U\       :  �J  �6   	         	  ���        ����
 � �����  �  @         ����   ( )          w � \`       [  �K  �C           	  ���        ����
 � �����  �  @         ����   * +          | � cd       |  &M  �P           	  ���        ����
 � �����  �  @         ����   , -          � � jh       �  RN  �]           	  ���       ����
 � �����  �  @         ����   . /          � � ql       �  ~O  jj           	  ���       ����
 � �����  �  @         ����   0 1          � � xp       �  �P  Nw           	  ���       ����
 � �����  �  @         ����   3 4          � � t        	  �Q  2�           	  ���       ����
 � �����  �  @         ����   5 6          � � �x       !	  S  �   ��       	  ���       ����
 � �����  �  @         ����   7 8          � � �|       B	  .T  ��   ��       	  ���       ����
 � �����  �  @         ����   9 :          � � ��       c	  ZU  ު   ��  	     	  ���       ����
 7  �  �  @         ����   * +          � � |j d     �
  
Z  x8            
  ���        ���� � �����  �  A         ����   , -          � � �o e     �
  T[  �G           
  ���        ���� � �����  �  A         ����   . /          � � �t f       �\  hW           
  ���        ���� � �����  �  A         ����   0 1          � � �y g     D  �]  �f           
  ���       ���� � �����  �  A         ����   2 3          � � �~ h     l  2_  Xv           
  ���       ���� � �����  �  A         ����   4 5          � � �� i     �  |`  Ѕ   ��       
  ���       ���� � �����  �  A         ����   7 8          � � �� j     �  �a  H�   ��       
  ���       ���� � �����  �  A         ����   9 :          � � �� k     �  c  ��   ��       
  ���       ���� � �����  �  A         ����   ; <          � � �� l     
  Zd  8�   ��       
  ���       ���� �����  �  A         ����   = >          � � �� m     2  �e  ��   ��  	     
  ���       ���� A  �  �  A         ����   . /          � � �� n     �  �j  \l              ���        ���� � �����  �  B         ����   0 1          � � �� o       4l  �~             ���        ���� � �����  �  B         ����   2 3          � � �� p     ?  �m  �             ���        ���� � �����  �  B         ����   4 5          � � �� q     n  o  4�   ��         ���       ���� � �����  �  B         ����   6 7          � � �� r     �  lp  |�   ��         ���       ���� � �����  �  B         ����   8 9          � �� s     �  �q  ��   ��         ���       ���� � �����  �  B         ����   ; <          � 	�� t     �  <s  �   ��         ���       ����  �����  �  B         ����   = >          � �� u     )  �t  T�   ��         ���       ���� �����  �  B         ����   ? @          � �� v     X  v  ��   ��         ���       ���� �����  �  B         ����   A B          � �� w     �  tw  �   ��  	       ���       ���� A  �  �  B         ����   2 3          � �� x     �  }  �              ���        ���� � �����  �  C         ����   4 5          � 	�� y     �  �~  l�              ���        ���� � �����  �  C         ����   6 7          � �� z     �   �  �   ��         ���        ���� � �����  �  C         ����   8 9          � �� {     &  ��     ��         ���       ���� � �����  �  C         ����   : ;          � �� |     ]  ,�  h,   ��         ���       ����  �����  �  C         ����   < =          � !�� }     �  ��  �A   ��         ���       ���� �����  �  C         ����   ? @          � '� ~     �  8�  W   ��         ���       ���� �����  �  C         ����   A B          � -	�        ��  dl   ��         ���       ���� �����  �  C         ����   C D          � 3� �     7  D�  ��   ��         ���       ���� �����  �  C         ����   E F          � 9� �     n  ʊ  �   ��  	       ���       ���� #K  �  �  C          ����                ! !            �  F       w        ���        ���� � ������������D          ����                ! &            �  �	       w       ���        ���� � ������������D          ����                ! +            �  �	       w       ���        ���� � ������������D          ����                ! 0            
  
       w       ���       ���� � ������������D          ����   	 
            ! 5            (  P
       w       ���       ���� � ������������D          ����                ! :            F  �
       w       ���       ���� � ������������D          ����                ! ?            d  �
       w       ���       ���� � ������������D          ����                ! D            �         w       ���       ���� � ������������D          ����                ! I            �  @       w       ���       ���� � ������������D          ����                ! N            �  |       w	       ���       ���� � ������������D          ����                $ <         /   6  �       x        ���        ���� � ������������E          ����                ' A         1   r  V       x       ���        ���� � ������������E          ����   	 
            * F         3   �  
       x       ���        ���� � ������������E          ����                - K         5   �  �       x       ���       ���� � ������������E          ����                0 P         6   &  r       x       ���       ���� � ������������E          ����                3 U         8   b  &       x       ���       ���� � ������������E          ����                6 Z         :   �  �       x       ���       ���� � ������������E          ����                9 _         <   �  �       x       ���       ���� � ������������E          ����                < d         >     B       x       ���       ���� � ������������E          ����                ? i         ?   R  �       x	       ���       ���� � ������������E          ����   	 
           + V         ^   B	  %       y        ���        ���� � ������������F         ����              ! / [         b   �	  p&       y       ���        ���� � ������������F         ����              $ 3 `         f   �	  �'       y       ���        ���� � ������������F         ����              ' 7 e         i   P
  @)       y       ���       ���� � ������������F         ����              * ; j         m   �
  �*       y       ���       ���� � ������������F         ����              - ? o         p     ,       y       ���       ���� � ������������F         ����              0 C t         t   ^  x-       y       ���       ���� � ������������F         ����              3 G y         x   �  �.       y       ���       ���� � ������������F         ����              6 K ~         {     H0       y       ���       ���� � ������������F         ����              9 O �            l  �1       y	       ���       ���� � ������������F          ����              & < o        �   �  $E       z        ���        ���� � ������������G         ����              ) @ u        �   L  |G       z       ���        ���� � ������������G         ����              , D {         �   �  �I       z       ���        ���� � ������������G         ����              / H � #       �   <  ,L       z       ���       ���� � ������������G         ����              2 L � &       �   �  �N       z       ���       ���� � ������������G         ����              5 P � )       �   ,  �P       z       ���       ���� � ������������G         ����              8 T � ,       �   �  4S       z       ���       ���� � ������������G         ����              ; X � /       �     �U       z       ���       ���� � ������������G         ����              > \ � 2       �   �  �W       z       ���       ���� � ������������G         ����     !          A ` � 5       �     <Z       z	       ���       ���� � ������������G          ����              - L � !       2  �  �w       {        ���        ���� � ������������H         ����              0 P � $       ;  �  {       {       ���        ���� � ������������H         ����              3 T � '       D    �~       {       ���        ���� � ������������H         ����              6 X � *       M  �  �       {       ���       ���� � ������������H         ����              9 \ � -       V  D  ��       {       ���       ���� � ������������H         ����              < ` � 0       _  �  �       {       ���       ���� � ������������H         ����              ? d � 3       h  p  ��       {       ���       ���� � ������������H         ����     !          B h � 6       q    $�       {       ���       ���� � ������������H         ����   " #          E l � 9       z  �  ��    
   {       ���       ���� � ������������H         ����   $ %          H p � <       �  2  ,�    	   {	       ���       ���� � ������������H          ����              4 [ � (       �  �  ��       |        ���        ���� � ������������I         ����              8 _ � +       �  >  ��       |       ���        ���� � ������������I         ����              < c � .         �  ��       |       ���        ���� � ������������I         ����              @ g � 1         �  ��       |       ���       ���� � ������������I         ����              D k � 4         Z  v�       |       ���       ���� � ������������I         ����     !          H o � 7       ,    b�       |       ���       ���� � ������������I         ����   " #          L s � :       9  �  N�       |       ���       ���� � ������������I         ����   $ %          P w � =       E  v   :�    	   |       ���       ���� � ������������I         ����   & '          T { � @       R  *!  &�       |       ���       ���� � ������������I         ����   ( )          X  � C       ^  �!  �       |	       ���       ���� � ������������I         ����              D j � .       �  �$  p%      }        ���        ���� � �����  �  J         ����              H o � 2          �%   ,      }       ���        ���� � �����  �  J         ����              L t � 6         R&  �2      }       ���        ���� � �����  �  J         ����               P y � :       !  $'   9      }       ���       ���� � �����  �  J         ����   ! "          T ~ � >       2  �'  �?      }       ���       ���� � �����  �  J         ����   $ %          X � � B       C  �(  @F   	   }       ���       ���� � �����  �  J         ����   & '          \ � � F       T  �)  �L      }       ���       ���� � �����  �  J         ����   ( )          ` � � J       d  l*  `S      }       ���       ���� � �����  �  J         ����   * +          d � N       u  >+  �Y      }       ���       ���� � �����  �  J         ����   , -          h � 
R       �  ,  �`      }	       ���       ���� � �����  �  J         ����              T � � >       B  X/  �      ~        ���        ���� � �����  �  K         ����               X � � B       X  H0  ��      ~       ���        ���� � �����  �  K         ����   ! "          \ � F       n  81  ��      ~       ���        ���� � �����  �  K         ����   # $          ` � 	J       �  (2  h�   	   ~       ���       ���� � �����  �  K         ����   % &          d � N       �  3  ��      ~       ���       ���� � �����  �  K         ����   ' (          h � R       �  4  H�      ~       ���       ���� � �����  �  K         ����   * +          l � V       �  �4  ��      ~       ���       ���� � �����  �  K         ����   , -          p � %Z       �  �5  (�      ~       ���       ���� � �����  �  K         ����   . /          t � ,^       �  �6  ��      ~       ���       ���� � �����  �  K         ����   0 1          x � 3b         �7  �      ~	       ���       ���� � -  �  �  K         ����   ! "          c � M       �  �;  PS            	  ���        ����	 � �����  �  L         ����   # $          g � $Q         �<  �]   
        	  ���        ����	 � �����  �  L         ����   % &          k � +U       *  �=  hh           	  ���        ����	 � �����  �  L         ����   ' (          o � 2Y       E  �>  �r           	  ���       ����	 � �����  �  L         ����   ) *          s � 9]       `  �?  �}           	  ���       ����	 � �����  �  L         ����   + ,          w � @a       {  �@  �           	  ���       ����	 � �����  �  L         ����   . /          { � Ge       �  �A  ��           	  ���       ����	 � �����  �  L         ����   0 1           � Ni       �  �B  $�           	  ���       ����	 � �����  �  L         ����   2 3          � � Um       �  �C  ��            	  ���       ����	 � �����  �  L         ����   4 5          � � \q       �  E  <�   ��  	     	  ���       ����	 � 7  �  �  L         ����   % &          r � E\         >I  �%   	   �      
  ���        ����
 � �����  �  M         ����   ' (          w � L`       /  jJ  �2      �     
  ���        ����
 � �����  �  M         ����   ) *          | � Sd       P  �K  r?      �     
  ���        ����
 � �����  �  M         ����   + ,          � � Zh       q  �L  VL      �     
  ���       ����
 � �����  �  M         ����   - .          � � al       �  �M  :Y      �     
  ���       ����
 � �����  �  M         ����   / 0          � � hp       �  O  f      �     
  ���       ����
 � �����  �  M         ����   2 3          � � ot       �  FP  s      �     
  ���       ����
 � �����  �  M         ����   4 5          � � vx       �  rQ  �   ��  �     
  ���       ����
 � �����  �  M         ����   6 7          � � }|       	  �R  ʌ   ��  �     
  ���       ����
 � �����  �  M         ����   8 9          � � ��       7	  �S  ��   ��  �	     
  ���       ����
 7  �  �  M         ����   ) *          � � lj d     �
  zX  �%      �        ���        ���� � �����  �  N         ����   + ,          � � so e     �
  �Y  05      �       ���        ���� � �����  �  N         ����   - .          � � zt f     �
  [  �D      �       ���        ���� � �����  �  N         ����   / 0          � � �y g       X\   T      �       ���       ���� � �����  �  N         ����   1 2          � � �~ h     <  �]  �c      �       ���       ���� � �����  �  N         ����   3 4          � � �� i     d  �^  s   ��  �       ���       ���� � �����  �  N         ����   6 7          � � �� j     �  6`  ��   ��  �       ���       ���� � �����  �  N         ����   8 9          � � �� k     �  �a   �   ��  �       ���       ���� � �����  �  N         ����   : ;          � � �� l     �  �b  x�   ��  �       ���       ���� �����  �  N         ����   < =          � � �� m       d  �   ��  �	       ���       ���� A  �  �  N         ����   - .          � � �� n     �  <i  X      �        ���        ���� � �����  �  O         ����   / 0          � � �� o     �  �j  Tj      �       ���        ���� � �����  �  O         ����   1 2          � � �� p       l  �|      �       ���        ���� � �����  �  O         ����   3 4          � � �� q     :  tm  �   ��  �       ���       ���� � �����  �  O         ����   5 6          � � �� r     i  �n  ,�   ��  �       ���       ���� � �����  �  O         ����   7 8          � �� s     �  Dp  t�   ��  �       ���       ���� � �����  �  O         ����   : ;          � 	�� t     �  �q  ��   ��  �       ���       ����  �����  �  O         ����   < =          � �� u     �  s  �   ��  �       ���       ���� �����  �  O         ����   > ?          � �� v     $  |t  L�   ��  �       ���       ���� �����  �  O         ����   @ A          � �� w     S  �u  ��   ��  �	       ���       ���� A  �  �  O         ����   1 2          � �� x     J  �{  8�      �        ���        ���� � �����  �  P         ����   3 4          � 	�� y     �  
}  ��       �       ���        ���� � �����  �  P         ����   5 6          � �� z     �  �~  ��   ��  �       ���        ���� � �����  �  P         ����   7 8          � �� {     �  �  4   ��  �       ���       ���� � �����  �  P         ����   9 :          � �� |     %  ��  �   ��  �       ���       ����  �����  �  P         ����   ; <          � !�� }     [  "�  �+   ��  �       ���       ���� �����  �  P         ����   > ?          � '�� ~     �  ��  0A   ��  �       ���       ���� �����  �  P         ����   @ A          � -��      �  .�  �V   ��  �       ���       ���� �����  �  P         ����   B C          � 3� �     �  ��  �k   ��  �       ���       ���� �����  �  P         ����   D E          � 9	� �     6  :�  ,�   ��  �	       ���       ���� #K  �  �  P          ����                - -         2   `	  �       �      �   �        ���� � ������������Q          ����                - 2         0   ~	  �       �     �   �        ���� � ������������Q          ����                - 7         1   �	  8       �     �   �        ���� � ������������Q          ����    	            - <         1   �	  t       �     �   �       ���� � ������������Q          ����   
             - A         2   �	  �       �     �   �       ���� � ������������Q          ����                - F         3   �	  �       �     �   �       ���� � ������������Q          ����                - K         3   
  (       �     �   �       ���� � ������������Q          ����                - P         4   2
  d       �     �   �       ���� � ������������Q          ����                - U         4   P
  �       �     �   �       ���� � ������������Q          ����                - Z         5   n
  �       �	     �   �       ���� � ������������Q          ����                $ H         S   �
  �        �      �   �        ���� � ������������R          ����    	            ' M         U   "  f!       �     �   �        ���� � ������������R          ����   
             * R         W   ^  "       �     �   �        ���� � ������������R          ����                - W         Y   �  �"       �     �   �       ���� � ������������R          ����                0 \         Z   �  �#       �     �   �       ���� � ������������R          ����                3 a         \     6$       �     �   �       ���� � ������������R          ����                6 f         ^   N  �$       �     �   �       ���� � ������������R          ����                9 k         `   �  �%       �     �   �       ���� � ������������R          ����                < p         b   �  R&       �     �   �       ���� � ������������R          ����                ? u         c     '       �	     �   �       ���� � ������������R         ����   
            + b         �   �  �7       �      �   �        ���� � ������������S         ����              ! / g         �   L  09       �     �   �        ���� � ������������S         ����              $ 3 l         �   �  �:       �     �   �        ���� � ������������S         ����              ' 7 q         �       <       �     �   �       ���� � ������������S         ����              * ; v         �   Z  h=       �     �   �       ���� � ������������S         ����              - ? {         �   �  �>       �     �   �       ���� � ������������S         ����              0 C �         �     8@       �     �   �       ���� � ������������S         ����              3 G �         �   h  �A       �     �   �       ���� � ������������S         ����              6 K �         �   �  C       �     �   �       ���� � ������������S         ����              9 O �         �     pD       �	     �   �       ���� � ������������S         ����              & < {        �   �  �\       �      �   �        ���� � ������������T         ����              ) @ �        �   �  �^       �     �   �        ���� � ������������T         ����              , D �         �   t  Da       �     �   �        ���� � ������������T         ����              / H � #       �   �  �c       �     �   �       ���� � ������������T         ����              2 L � &         d  �e       �     �   �       ���� � ������������T         ����              5 P � )         �  Lh       �     �   �       ���� � ������������T         ����              8 T � ,         T  �j       �     �   �       ���� � ������������T         ����              ; X � /         �  �l       �     �   �       ���� � ������������T         ����               > \ � 2         D  To       �     �   �       ���� � ������������T         ����   ! "          A ` � 5       #  �  �q       �	     �   �       ���� � ������������T         ����              - L � !       z  �  ��       �      �   �        ���� � ������������U         ����              0 P � $       �  2  ,�       �     �   �        ���� � ������������U         ����              3 T � '       �  �  ��       �     �   �        ���� � ������������U         ����              6 X � *       �  ^  4�       �     �   �       ���� � ������������U         ����              9 \ � -       �  �  ��       �     �   �       ���� � ������������U         ����              < ` � 0       �  �  <�       �     �   �       ���� � ������������U         ����               ? d � 3       �     ��       �     �   �       ���� � ������������U         ����   ! "          B h � 6       �  �  D�       �     �   �       ���� � ������������U         ����   # $          E l � 9       �  L  ȯ    
   �     �   �       ���� � ������������U         ����   % &          H p � <       �  �  L�    	   �	     �   �       ���� � ������������U         ����              4 [ � (       A  :   ��       �      �   �        ���� � ������������V         ����              8 _ � +       N  �   ��       �     �   �        ���� � ������������V         ����              < c � .       Z  �!  n�       �     �   �        ���� � ������������V         ����              @ g � 1       g  V"  Z�       �     �   �       ���� � ������������V         ����              D k � 4       s  
#  F�       �     �   �       ���� � ������������V         ����   ! "          H o � 7       �  �#  2�       �     �   �       ���� � ������������V         ����   # $          L s � :       �  r$  �       �     �   �       ���� � ������������V         ����   % &          P w � =       �  &%  
   	   �     �   �       ���� � ������������V         ����   ' (          T { � @       �  �%  �      �     �   �       ���� � ������������V         ����   ) *          X  � C       �  �&  �      �	     �   �       ���� � ������������V         ����              D j � .       O  ^)  �J      �      �   �        ���� � �����  �  W         ����              H o � 2       `  0*  �Q      �     �   �        ���� � �����  �  W         ����              L t � 6       p  +  X      �     �   �        ���� � �����  �  W         ����     !          P y � :       �  �+  �^      �     �   �       ���� � �����  �  W         ����   " #          T ~ � >       �  �,  0e      �     �   �       ���� � �����  �  W         ����   $ %          X � � B       �  x-  �k   	   �     �   �       ���� � �����  �  W         ����   ' (          \ � F       �  J.  Pr      �     �   �       ���� � �����  �  W         ����   ) *          ` � 
J       �  /  �x      �     �   �       ���� � �����  �  W         ����   + ,          d � N       �  �/  p      �     �   �       ���� � �����  �  W         ����   - .          h � R       �  �0   �      �	     �   �       ���� � �����  �  W         ����              T �  >       �  4  H�      �      �   �        ���� � �����  �  X         ����     !          X � B       �  �4  ��      �     �   �        ���� � �����  �  X         ����   " #          \ � F       �  �5  (�      �     �   �        ���� � �����  �  X         ����   $ %          ` � J       �  �6  ��   	   �     �   �       ���� � �����  �  X         ����   & '          d � N         �7  �      �     �   �       ���� � �����  �  X         ����   ( )          h � #R         �8  x�      �     �   �       ���� � �����  �  X         ����   + ,          l � *V       0  �9  �      �     �   �       ���� � �����  �  X         ����   - .          p � 1Z       F  �:  X      �     �   �       ���� � �����  �  X         ����   / 0          t � 8^       [  �;  �      �     �   �       ���� � �����  �  X         ����   1 2          x � ?b       q  x<  8       �	     �   �       ���� � -  �  �  X         ����   " #          c � )M       l  8@  0�      �      �   �        ����	 � �����  �  Y         ����   $ %          g � 0Q       �  FA  ��   
   �     �   �        ����	 � �����  �  Y         ����   & '          k � 7U       �  TB  H�      �     �   �        ����	 � �����  �  Y         ����   ( )          o � >Y       �  bC  ԡ      �     �   �       ����	 � �����  �  Y         ����   * +          s � E]       �  pD  `�      �     �   �       ����	 � �����  �  Y         ����   , -          w � La       �  ~E  �      �     �   �       ����	 � �����  �  Y         ����   / 0          { � Se         �F  x�      �     �   �       ����	 � �����  �  Y         ����   1 2           � Zi       )  �G  �      �     �   �       ����	 � �����  �  Y         ����   3 4          � � am       D  �H  ��       �     �   �       ����	 � �����  �  Y         ����   5 6          � � hq       _  �I  �   ��  �	     �   �       ����	 � 7  �  �  Y         ����   & '          r � Q\       �  �M  :Y   	   �      �   �        ����
 � �����  �  Z         ����   ( )          w � X`       �  O  f      �     �   �        ����
 � �����  �  Z         ����   * +          | � _d       �  FP  s      �     �   �        ����
 � �����  �  Z         ����   , -          � � fh       �  rQ  �      �     �   �       ����
 � �����  �  Z         ����   . /          � � ml       	  �R  ʌ      �     �   �       ����
 � �����  �  Z         ����   0 1          � � tp       7	  �S  ��      �     �   �       ����
 � �����  �  Z         ����   3 4          � � {t       X	  �T  ��      �     �   �       ����
 � �����  �  Z         ����   5 6          � � �x       y	  "V  v�   ��  �     �   �       ����
 � �����  �  Z         ����   7 8          � � �|       �	  NW  Z�   ��  �     �   �       ����
 � �����  �  Z         ����   9 :          � � ��       �	  zX  >�   ��  �	     �   �       ����
 7  �  �  Z         ����   * +          � � xj d     .  *]  �]      �      �   �        ���� � �����  �  [         ����   , -          � � o e     U  t^  pm      �     �   �        ���� � �����  �  [         ����   . /          � � �t f     }  �_  �|      �     �   �        ���� � �����  �  [         ����   0 1          � � �y g     �  a  `�      �     �   �       ���� � �����  �  [         ����   2 3          � � �~ h     �  Rb  ؛      �     �   �       ���� � �����  �  [         ����   4 5          � � �� i     �  �c  P�   ��  �     �   �       ���� � �����  �  [         ����   7 8          � � �� j       �d  Ⱥ   ��  �     �   �       ���� � �����  �  [         ����   9 :          � � �� k     C  0f  @�   ��  �     �   �       ���� � �����  �  [         ����   ; <          � � �� l     j  zg  ��   ��  �     �   �       ���� �����  �  [         ����   = >          � � �� m     �  �h  0�   ��  �	     �   �       ���� A  �  �  [         ����   . /          � � �� n     J  �m  ��      �      �   �        ���� � �����  �  \         ����   0 1          � � �� o     y  To  D�      �     �   �        ���� � �����  �  \         ����   2 3          � � �� p     �  �p  ��      �     �   �        ���� � �����  �  \         ����   4 5          � � �� q     �  $r  ��   ��  �     �   �       ���� � �����  �  \         ����   6 7          � � �� r       �s  �   ��  �     �   �       ���� � �����  �  \         ����   8 9          � �� s     4  �t  d�   ��  �     �   �       ���� � �����  �  \         ����   ; <          � 	�� t     c  \v  �   ��  �     �   �       ����  �����  �  \         ����   = >          � �� u     �  �w  �   ��  �     �   �       ���� �����  �  \         ����   ? @          � �� v     �  ,y  <'   ��  �     �   �       ���� �����  �  \         ����   A B          � �� w     �  �z  �9   ��  �	     �   �       ���� A  �  �  \         ����   2 3          � �� x     �  4�  �      �      �   �        ���� � �����  �  ]         ����   4 5          � 	�� y     )  ��  ,       �     �   �        ���� � �����  �  ]         ����   6 7          � �� z     `  @�  �-   ��  �     �   �        ���� � �����  �  ]         ����   8 9          � �� {     �  Ƅ  �B   ��  �     �   �       ���� � �����  �  ]         ����   : ;          � �� |     �  L�  (X   ��  �     �   �       ����  �����  �  ]         ����   < =          � !�� }       ҇  |m   ��  �     �   �       ���� �����  �  ]         ����   ? @          � '�� ~     :  X�  Ђ   ��  �     �   �       ���� �����  �  ]         ����   A B          � -�      q  ފ  $�   ��  �     �   �       ���� �����  �  ]         ����   C D          � 3� �     �  d�  x�   ��  �     �   �       ���� �����  �  ]         ����   E F          � 9� �     �  �  ��   ��  �	     �   �       ���� #K  �  �  ]            ��                 @ @        �����
  �               � !   �        ���� � ������������^            ��                 @ E        ����               � !   �        ���� � ������������^            ��                 @ J        ����,  X             � !   �        ���� � ������������^            ��    	             @ O        ����J  �             � !   �        ���� � ������������^            ��   
              @ T        ����h  �             � !   �        ���� � ������������^            ��                 @ Y        �����               � !   �        ���� � ������������^            ��                 @ ^        �����  H             � !   �        ���� � ������������^            ��                 @ c        �����  �             � !   �        ���� � ������������^            ��                 @ h        �����  �             � !   �        ���� � ������������^            ��                 @ m        �����  �        	     � !   �        ���� � ������������^           ��                 $ [   (     ����v  b%              � !   �        ���� � ������������_           ��    	             ' `   (     �����  &             � !   �        ���� � ������������_           ��   
              * e   (     �����  �&             � !   �        ���� � ������������_           ��                 - j   (     ����*  ~'             � !   �        ���� � ������������_           ��                 0 o   (     ����f  2(             � !   �        ���� � ������������_           ��                 3 t   (     �����  �(             � !   �        ���� � ������������_           ��                 6 y   (     �����  �)             � !   �        ���� � ������������_           ��                 9 ~   (     ����  N*             � !   �        ���� � ������������_           ��                 < �   (     ����V  +             � !   �        ���� � ������������_           ��                 ? �   (     �����  �+        	     � !   �        ���� � ������������_          ��   
             + u   2     �����  >        	      � !   �        ���� � ������������`          ��               ! / z   2     �����  p?        	     � !   �        ���� � ������������`          ��               $ 3    2     ����6  �@        	     � !   �        ���� � ������������`          ��               ' 7 �   2     �����  @B        	     � !   �        ���� � ������������`          ��               * ; �   2     �����  �C        	     � !   �        ���� � ������������`          ��               - ? �   2     ����D  E        	     � !   �        ���� � ������������`          ��               0 C �   2     �����  xF        	     � !   �        ���� � ������������`          ��               3 G �   2     �����  �G        	     � !   �        ���� � ������������`          ��               6 K �   2     ����R  HI        	     � !   �        ���� � ������������`          ��               9 O �   2     �����  �J        		     � !   �        ���� � ������������`         	 ��               & < �  <     ����  dd        
      � !   �        ���� � ������������a         	 ��               ) @ �  <     �����  �f        
     � !   �        ���� � ������������a         	 ��               , D �   <     ����  i        
     � !   �        ���� � ������������a         	 ��               / H � # <     ����|  lk        
     � !   �        ���� � ������������a         	 ��               2 L � & <     �����  �m        
     � !   �        ���� � ������������a         	 ��               5 P � ) <     ����l  p        
     � !   �        ���� � ������������a         	 ��               8 T � , <     �����  tr        
     � !   �        ���� � ������������a         	 ��               ; X � / <     ����\  �t        
     � !   �        ���� � ������������a         	 ��                > \ � 2 <     �����  $w        
     � !   �        ���� � ������������a         	 ��   ! "           A ` � 5 <     ����L  |y        
	     � !   �        ���� � ������������a         
 ��               - L � ! F     ����,  �              � !   �        ���� � ������������b         
 ��               0 P � $ F     �����  ��             � !   �        ���� � ������������b         
 ��               3 T � ' F     ����X  �             � !   �        ���� � ������������b          ��               6 X � * F     �����  ��             � !   �        ���� � ������������b          ��               9 \ � - F     �����  �             � !   �        ���� � ������������b          ��               < ` � 0 F     ����  ��             � !   �        ���� � ������������b          ��                ? d � 3 F     �����   �             � !   �        ���� � ������������b          ��   ! "           B h � 6 F     ����F  ��             � !   �        ���� � ������������b          ��   # $           E l � 9 F     �����  (�             � !   �        ���� � ������������b          ��   % &           H p � < F     ����r  ��        	     � !   �        ���� � ������������b          ��               4 [ � ( P     �����!  ��              � !   �        ���� � ������������c          ��               8 _ � + P     ����~"  r�             � !   �        ���� � ������������c          ��               < c � . P     ����2#  ^�             � !   �        ���� � ������������c          ��               @ g � 1 P     �����#  J�             � !   �        ���� � ������������c          ��               D k � 4 P     �����$  6             � !   �        ���� � ������������c          ��   ! "           H o � 7 P     ����N%  "            � !   �        ���� � ������������c          ��   # $           L s � : P     ����&  
            � !   �        ���� � ������������c          ��   % &           P w � = P     �����&  �            � !   �        ���� � ������������c          ��   ' (           T { @ P     ����j'  �            � !   �        ���� � ������������c          ��   ) *           X  C P     ����(  �       	     � !   �        ���� � ������������c          ��               D j � . Z     �����*  pW             � !   �        ���� � �����  �  d          ��               H o � 2 Z     �����+   ^            � !   �        ���� � �����  �  d          ��               L t � 6 Z     �����,  �d            � !   �        ���� � �����  �  d          ��     !           P y : Z     ����d-   k            � !   �        ���� � �����  �  d          ��   " #           T ~ > Z     ����6.  �q            � !   �        ���� � �����  �  d          ��   $ %           X � B Z     ����/  @x            � !   �        ���� � �����  �  d          ��   ' (           \ � F Z     �����/  �~            � !   �        ���� � �����  �  d          ��   ) *           ` � J Z     �����0  `�            � !   �        ���� � �����  �  d          ��   + ,           d � #N Z     ����~1  ��            � !   �        ���� � �����  �  d          ��   - .           h � )R Z     ����P2  ��       	     � !   �        ���� � �����  �  d          ��               T � > d     �����5  X�             � !   �        ���� � �����  �  e          ��     !           X � B d     �����6  ��            � !   �        ���� � �����  �  e          ��   " #           \ � !F d     ����x7  8�            � !   �        ���� � �����  �  e          ��   $ %           ` � (J d     ����h8  ��            � !   �        ���� � �����  �  e          ��   & '           d � /N d     ����X9              � !   �        ���� � �����  �  e          ��   ( )           h � 6R d     ����H:  �            � !   �        ���� � �����  �  e          ��   + ,           l � =V d     ����8;  �            � !   �        ���� � �����  �  e          ��   - .           p � DZ d     ����(<  h            � !   �        ���� � �����  �  e          ��   / 0           t � K^ d     ����=  �%            � !   �        ���� � �����  �  e          ��   1 2           x � Rb d     ����>  H.       	     � !   �        ���� � �����  �  e          ��   " #           c � <M n     �����A  Б             � !   �        ����	 � �����  �  f          ��   $ %           g � CQ n     �����B  \�            � !   �        ����	 � �����  �  f          ��   & '           k � JU n     �����C  �            � !   �        ����	 � �����  �  f          ��   ( )           o � QY n     �����D  t�            � !   �        ����	 � �����  �  f          ��   * +           s � X] n     ���� F   �            � !   �        ����	 � �����  �  f          ��   , -           w � _a n     ����G  ��            � !   �        ����	 � �����  �  f          ��   / 0           { � fe n     ����H  �            � !   �        ����	 � �����  �  f          ��   1 2            � mi n     ����*I  ��            � !   �        ����	 � �����  �  f          ��   3 4           � � tm n     ����8J  0�            � !   �        ����	 � �����  �  f          ��   5 6           � � {q n     ����FK  ��       	     � !   �        ����	 � �����  �  f          ��   & '           r � d\ x     ����~O  jj             � !   �        ����
 � �����  �  g          ��   ( )           w � k` x     �����P  Nw            � !   �        ����
 � �����  �  g          ��   * +           | � rd x     �����Q  2�            � !   �        ����
 � �����  �  g          ��   , -           � � yh x     ����S  �            � !   �        ����
 � �����  �  g          ��   . /           � � �l x     ����.T  ��            � !   �        ����
 � �����  �  g          ��   0 1           � � �p x     ����ZU  ު            � !   �        ����
 � �����  �  g          ��   3 4           � � �t x     �����V  ·            � !   �        ����
 � �����  �  g          ��   5 6           � � �x x     �����W  ��            � !   �        ����
 � �����  �  g          ��   7 8           � � �| x     �����X  ��            � !   �        ����
 � �����  �  g          ��   9 :           � � �� x     ����
Z  n�       	     � !   �        ����
 �����  �  g          ��   * +           � � �j �     �����^  �p             � !   �        ���� � �����  �  h          ��   , -           � � �o �     ����`  0�            � !   �        ���� � �����  �  h          ��   . /           � � �t �     ����Na  ��            � !   �        ���� � �����  �  h          ��   0 1           � � �y �     �����b   �            � !   �        ���� � �����  �  h          ��   2 3           � � �~ �     �����c  ��            � !   �        ���� � �����  �  h          ��   4 5           � � �� �     ����,e  �            � !   �        ���� � �����  �  h          ��   7 8           � � �� �     ����vf  ��            � !   �        ���� � �����  �  h          ��   9 :           � � �� �     �����g   �            � !   �        ���� � �����  �  h          ��   ; <           � � �� �     ����
i  x�            � !   �        ���� �����  �  h          ��   = >           � � �� �     ����Tj  ��       	     � !   �        ���� �����  �  h           ��   . /           � � �� �     ����|o  L�             � !   �        ���� � �����  �  i           ��   0 1           � � �� �     �����p  ��            � !   �        ���� � �����  �  i           ��   2 3           � � �� �     ����Lr  ��            � !   �        ���� � �����  �  i         ! ��   4 5           � � �� �     �����s  $�            � !   �        ���� � �����  �  i         ! ��   6 7           � � �� �     ����u  l�            � !   �        ���� � �����  �  i         ! ��   8 9           � �� �     �����v  �            � !   �        ���� � �����  �  i         " ��   ; <           � 	�� �     �����w  �            � !   �        ����  �����  �  i         " ��   = >           � �� �     ����Ty  D)            � !   �        ���� �����  �  i         " ��   ? @           � �� �     �����z  �;            � !   �        ���� �����  �  i         # ��   A B           � �� �     ����$|  �M       	     � !   �        ���� �����  �  i         $ ��   2 3           � �� �     ����ā  �             � !   �        ���� � �����  �  j         $ ��   4 5           � 	�� �     ����J�  .            � !   �        ���� � �����  �  j         $ ��   6 7           � �� �     ����Є  `C            � !   �        ���� � �����  �  j         $ ��   8 9           � �� �     ����V�  �X            � !   �        ���� � �����  �  j         $ ��   : ;           �  � �     ����܇  n            � !   �        ����  �����  �  j         $ ��   < =           � !� �     ����b�  \�            � !   �        ���� �����  �  j         $ ��   ? @           � '� �     �����  ��            � !   �        ���� �����  �  j         $ ��   A B           � -� �     ����n�  �            � !   �        ���� �����  �  j         $ ��   C D           � 3 � �     �����  X�            � !   �        ���� �����  �  j         $ ��   E F           � 9(� �     ����z�  ��       	     � !   �        ���� #�����  �  j          ����	                           ����  .J       (      ��! ���        ���� � ������������k          ����	                  $         ����.  \       (     ��! ���        ���� � ������������k          ����	                  )         ����L  �       (     ��! ���        ���� � ������������k          ����	                  .         ����j  �       (     ��! ���       ���� � ������������k          ����	   	 
              3         �����         (     ��! ���       ���� � ������������k          ����	                  8         �����  L       (     ��! ���       ���� � ������������k          ����	                  =         �����  �       (     ��! ���       ���� � ������������k          ����	                  B         �����  �       (     ��! ���       ���� � ������������k          ����	                  G         ����           (     ��! ���       ���� � ������������k          ����	                  L         ����  <       (	     ��! ���       ���� � ������������k          ����	                 $ :         �����  �.       )      ��! ���        ���� � ������������l          ����	                 ' ?         �����  v/       )     ��! ���        ���� � ������������l          ����	   	 
             * D         ����  *0       )     ��! ���        ���� � ������������l          ����	                 - I         ����J  �0       )     ��! ���       ���� � ������������l          ����	                 0 N         �����  �1       )     ��! ���       ���� � ������������l          ����	                 3 S         �����  F2       )     ��! ���       ���� � ������������l          ����	                 6 X         �����  �2       )     ��! ���       ���� � ������������l          ����	                 9 ]         ����:  �3       )     ��! ���       ���� � ������������l          ����	                 < b         ����v  b4       )     ��! ���       ���� � ������������l          ����	                 ? g         �����  5       )	     ��! ���       ���� � ������������l         ����	   	 
            + T         �����  �J       *      ��! ���        ���� � ������������m         ����	               ! / Y         �����  �K       *     ��! ���        ���� � ������������m         ����	               $ 3 ^         ����V  XM       *     ��! ���        ���� � ������������m         ����	               ' 7 c         �����  �N       *     ��! ���       ���� � ������������m         ����	               * ; h         ����
  (P       *     ��! ���       ���� � ������������m         ����	               - ? m         ����d  �Q       *     ��! ���       ���� � ������������m         ����	               0 C r         �����  �R       *     ��! ���       ���� � ������������m         ����	               3 G w         ����  `T       *     ��! ���       ���� � ������������m         ����	               6 K |         ����r  �U       *     ��! ���       ���� � ������������m         ����	               9 O �         �����  0W       *	     ��! ���       ���� � ������������m         ����	               & < m        ����4  t       +      ��! ���        ���� � ������������n         ����	               ) @ s        �����  \v       +     ��! ���        ���� � ������������n         ����	               , D y         ����$  �x       +     ��! ���        ���� � ������������n         ����	               / H  #       �����  {       +     ��! ���       ���� � ������������n         ����	               2 L � &       ����  d}       +     ��! ���       ���� � ������������n         ����	               5 P � )       �����  �       +     ��! ���       ���� � ������������n         ����	               8 T � ,       ����  �       +     ��! ���       ���� � ������������n         ����	               ; X � /       ����|  l�       +     ��! ���       ���� � ������������n         ����	               > \ � 2       �����  Ć       +     ��! ���       ���� � ������������n         ����	     !           A ` � 5       ����l  �       +	     ��! ���       ���� � ������������n         ����	               - L � !       ����L  ȯ       ,      ��! ���        ���� � ������������o         ����	               0 P � $       �����  L�       ,     ��! ���        ���� � ������������o         ����	               3 T � '       ����x  ж       ,     ��! ���        ���� � ������������o         ����	               6 X � *       ����  T�       ,     ��! ���       ���� � ������������o         ����	               9 \ � -       �����  ؽ       ,     ��! ���       ���� � ������������o         ����	               < ` � 0       ����:   \�       ,     ��! ���       ���� � ������������o         ����	               ? d � 3       �����   ��       ,     ��! ���       ���� � ������������o         ����	     !           B h � 6       ����f!  d�       ,     ��! ���       ���� � ������������o         ����	   " #           E l � 9       �����!  ��    
   ,     ��! ���       ���� � ������������o         ����	   $ %           H p � <       �����"  l�    	   ,	     ��! ���       ���� � ������������o         ����	               4 [ � (       �����$  f      -      ��! ���        ���� � ������������p         ����	               8 _ � +       �����%  R      -     ��! ���        ���� � ������������p         ����	               < c � .       ����R&  >      -     ��! ���        ���� � ������������p         ����	               @ g � 1       ����'  *      -     ��! ���       ���� � ������������p         ����	               D k � 4       �����'        -     ��! ���       ���� � ������������p         ����	     !           H o � 7       ����n(        -     ��! ���       ���� � ������������p         ����	   " #           L s � :       ����")  �      -     ��! ���       ���� � ������������p         ����	   $ %           P w � =       �����)  �$   	   -     ��! ���       ���� � ������������p         ����	   & '           T { � @       �����*  �)      -     ��! ���       ���� � ������������p         ����	   ( )           X  � C       ����>+  �.      -	     ��! ���       ���� � ������������p         ����	               D j � .       ����.  pp      .      ��! ���        ���� � �����  �  q         ����	               H o � 2       �����.   w      .     ��! ���        ���� � �����  �  q         ����	               L t � 6       �����/  �}      .     ��! ���        ���� � �����  �  q         ����	                P y � :       �����0   �      .     ��! ���       ���� � �����  �  q         ����	   ! "           T ~ � >       ����V1  ��      .     ��! ���       ���� � �����  �  q         ����	   $ %           X � � B       ����(2  @�   	   .     ��! ���       ���� � �����  �  q         ����	   & '           \ � � F       �����2  З      .     ��! ���       ���� � �����  �  q         ����	   ( )           ` � � J       �����3  `�      .     ��! ���       ���� � �����  �  q         ����	   * +           d � N       �����4  �      .     ��! ���       ���� � �����  �  q         ����	   , -           h � R       ����p5  ��      .	     ��! ���       ���� � �����  �  q         ����	               T � � >       �����8  x�      /      ��! ���        ���� � �����  �  r         ����	                X � � B       �����9  �      /     ��! ���        ���� � �����  �  r         ����	   ! "           \ �  F       �����:  X      /     ��! ���        ���� � �����  �  r         ����	   # $           ` � J       �����;  �   	   /     ��! ���       ���� � �����  �  r         ����	   % &           d � N       ����x<  8       /     ��! ���       ���� � �����  �  r         ����	   ' (           h � R       ����h=  �(      /     ��! ���       ���� � �����  �  r         ����	   * +           l � V       ����X>  1      /     ��! ���       ���� � �����  �  r         ����	   , -           p � #Z       ����H?  �9      /     ��! ���       ���� � �����  �  r         ����	   . /           t � *^       ����8@  �A      /     ��! ���       ���� � �����  �  r         ����	   0 1           x � 1b       ����(A  hJ      /	     ��! ���       ���� � �����  �  r         ����	   ! "           c � M       �����D  �      0      ��! ���        ����	 � �����  �  s         ����	   # $           g � "Q       �����E  ��   
   0     ��! ���        ����	 � �����  �  s         ����	   % &           k � )U       ����G  (�      0     ��! ���        ����	 � �����  �  s         ����	   ' (           o � 0Y       ����H  ��      0     ��! ���       ����	 � �����  �  s         ����	   ) *           s � 7]       ���� I  @�      0     ��! ���       ����	 � �����  �  s         ����	   + ,           w � >a       ����.J  ��      0     ��! ���       ����	 � �����  �  s         ����	   . /           { � Ee       ����<K  X�      0     ��! ���       ����	 � �����  �  s         ����	   0 1            � Li       ����JL  ��      0     ��! ���       ����	 � �����  �  s         ����	   2 3           � � Sm       ����XM  p       0     ��! ���       ����	 � �����  �  s         ����	   4 5           � � Zq       ����fN  �   ��  0	     ��! ���       ����	 � �����  �  s         ����	   % &           r � C\       �����R  ʌ   	   1      ��! ���        ����
 � �����  �  t         ����	   ' (           w � J`       �����S  ��      1     ��! ���        ����
 � �����  �  t         ����	   ) *           | � Qd       �����T  ��      1     ��! ���        ����
 � �����  �  t         ����	   + ,           � � Xh       ����"V  v�      1     ��! ���       ����
 � �����  �  t         ����	   - .           � � _l       ����NW  Z�      1     ��! ���       ����
 � �����  �  t         ����	   / 0           � � fp       ����zX  >�      1     ��! ���       ����
 � �����  �  t         ����	   2 3           � � mt       �����Y  "�      1     ��! ���       ����
 � �����  �  t         ����	   4 5           � � tx       �����Z  �   ��  1     ��! ���       ����
 � �����  �  t         ����	   6 7           � � {|       �����[  ��   ��  1     ��! ���       ����
 � �����  �  t         ����	   8 9           � � ��       ����*]  �    ��  1	     ��! ���       ����
 �����  �  t         ����	   ) *           � � jj d     �����a  8�      2      ��! ���        ���� � �����  �  u         ����	   + ,           � � qo e     ����$c  ��      2     ��! ���        ���� � �����  �  u         ����	   - .           � � xt f     ����nd  (�      2     ��! ���        ���� � �����  �  u         ����	   / 0           � � y g     �����e  ��      2     ��! ���       ���� � �����  �  u         ����	   1 2           � � �~ h     ����g  �      2     ��! ���       ���� � �����  �  u         ����	   3 4           � � �� i     ����Lh  ��   ��  2     ��! ���       ���� � �����  �  u         ����	   6 7           � � �� j     �����i  �   ��  2     ��! ���       ���� � �����  �  u         ����	   8 9           � � �� k     �����j  �   ��  2     ��! ���       ���� � �����  �  u         ����	   : ;           � � �� l     ����*l  �   ��  2     ��! ���       ���� �����  �  u         ����	   < =           � � �� m     ����tm  p!   ��  2	     ��! ���       ���� �����  �  u         ����	   - .           � � �� n     �����r  ��      3      ��! ���        ���� � �����  �  v         ����	   / 0           � � �� o     ����t  4�      3     ��! ���        ���� � �����  �  v         ����	   1 2           � � �� p     ����lu  |�      3     ��! ���        ���� � �����  �  v         ����	   3 4           � � �� q     �����v  �   ��  3     ��! ���       ���� � �����  �  v         ����	   5 6           � � �� r     ����<x     ��  3     ��! ���       ���� � �����  �  v         ����	   7 8           � �� s     �����y  T-   ��  3     ��! ���       ���� � �����  �  v         ����	   : ;           � 	�� t     ����{  �?   ��  3     ��! ���       ����  �����  �  v         ����	   < =           � �� u     ����t|  �Q   ��  3     ��! ���       ���� �����  �  v         ����	   > ?           � �� v     �����}  ,d   ��  3     ��! ���       ���� �����  �  v         ����	   @ A           � �� w     ����D  tv   ��  3	     ��! ���       ���� �����  �  v         ����	   1 2           � �� x     �����  xD      4      ��! ���        ���� � �����  �  w         ����	   3 4           � 	�� y     ����j�  �Y       4     ��! ���        ���� � �����  �  w         ����	   5 6           � �� z     ������   o   ��  4     ��! ���        ���� � �����  �  w         ����	   7 8           � �� {     ����v�  t�   ��  4     ��! ���       ���� � �����  �  w         ����	   9 :           � �� |     ������  ș   ��  4     ��! ���       ����  �����  �  w         ����	   ; <           � !�� }     ������  �   ��  4     ��! ���       ���� �����  �  w         ����	   > ?           � '�� ~     �����  p�   ��  4     ��! ���       ���� �����  �  w         ����	   @ A           � -��      ������  ��   ��  4     ��! ���       ���� �����  �  w         ����	   B C           � 3�� �     �����  �   ��  4     ��! ���       ���� �����  �  w         ����	   D E           � 9� �     ������  l   ��  4	     ��! ���       ���� #�����  �  w          ����
                 ' '         �����  t1       �      ��! ���        ���� � ������������x          ����
                 ' ,         �����  <       �     ��! ���        ���� � ������������x          ����
                 ' 1         �����  x       �     ��! ���        ���� � ������������x          ����
                 ' 6         �����  �       �     ��! ���       ���� � ������������x          ����
   	 
             ' ;         �����  �       �     ��! ���       ���� � ������������x          ����
                 ' @         ����  ,       �     ��! ���       ���� � ������������x          ����
                 ' E         ����4  h       �     ��! ���       ���� � ������������x          ����
                 ' J         ����R  �       �     ��! ���       ���� � ������������x          ����
                 ' O         ����p  �       �     ��! ���       ���� � ������������x          ����
                 ' T         �����         �	     ��! ���       ���� � ������������x          ����
                 $ B         ����  *       �      ��! ���        ���� � ������������y          ����
                 ' G         ����B  �*       �     ��! ���        ���� � ������������y          ����
   	 
             * L         ����~  z+       �     ��! ���        ���� � ������������y          ����
                 - Q         �����  .,       �     ��! ���       ���� � ������������y          ����
                 0 V         �����  �,       �     ��! ���       ���� � ������������y          ����
                 3 [         ����2  �-       �     ��! ���       ���� � ������������y          ����
                 6 `         ����n  J.       �     ��! ���       ���� � ������������y          ����
                 9 e         �����  �.       �     ��! ���       ���� � ������������y          ����
                 < j         �����  �/       �     ��! ���       ���� � ������������y          ����
                 ? o         ����"  f0       �	     ��! ���       ���� � ������������y         ����
   	 
            + \         ����  HD       �      ��! ���        ���� � ������������z         ����
               ! / a         ����l  �E       �     ��! ���        ���� � ������������z         ����
               $ 3 f         �����  G       �     ��! ���        ���� � ������������z         ����
               ' 7 k         ����   �H       �     ��! ���       ���� � ������������z         ����
               * ; p         ����z  �I       �     ��! ���       ���� � ������������z         ����
               - ? u         �����  PK       �     ��! ���       ���� � ������������z         ����
               0 C z         ����.  �L       �     ��! ���       ���� � ������������z         ����
               3 G          �����   N       �     ��! ���       ���� � ������������z         ����
               6 K �         �����  �O       �     ��! ���       ���� � ������������z         ����
               9 O �         ����<  �P       �	     ��! ���       ���� � ������������z         ����
               & < u        �����  4l       �      ��! ���        ���� � ������������{         ����
               ) @ {        ����  �n       �     ��! ���        ���� � ������������{         ����
               , D �         �����  �p       �     ��! ���        ���� � ������������{         ����
               / H � #       ����  <s       �     ��! ���       ���� � ������������{         ����
               2 L � &       �����  �u       �     ��! ���       ���� � ������������{         ����
               5 P � )       �����  �w       �     ��! ���       ���� � ������������{         ����
               8 T � ,       ����t  Dz       �     ��! ���       ���� � ������������{         ����
               ; X � /       �����  �|       �     ��! ���       ���� � ������������{         ����
               > \ � 2       ����d  �~       �     ��! ���       ���� � ������������{         ����
     !           A ` � 5       �����  L�       �	     ��! ���       ���� � ������������{         ����
               - L � !       �����  h�       �      ��! ���        ���� � ������������|         ����
               0 P � $       ����R  �       �     ��! ���        ���� � ������������|         ����
               3 T � '       �����  p�       �     ��! ���        ���� � ������������|         ����
               6 X � *       ����~  ��       �     ��! ���       ���� � ������������|         ����
               9 \ � -       ����  x�       �     ��! ���       ���� � ������������|         ����
               < ` � 0       �����  ��       �     ��! ���       ���� � ������������|         ����
               ? d � 3       ����@  ��       �     ��! ���       ���� � ������������|         ����
     !           B h � 6       �����  �       �     ��! ���       ���� � ������������|         ����
   " #           E l � 9       ����l   ��    
   �     ��! ���       ���� � ������������|         ����
   $ %           H p � <       ����!  �    	   �	     ��! ���       ���� � ������������|         ����
               4 [ � (       ����Z#  v�       �      ��! ���        ���� � ������������}         ����
               8 _ � +       ����$  b�       �     ��! ���        ���� � ������������}         ����
               < c � .       �����$  N      �     ��! ���        ���� � ������������}         ����
               @ g � 1       ����v%  :      �     ��! ���       ���� � ������������}         ����
               D k � 4       ����*&  &      �     ��! ���       ���� � ������������}         ����
     !           H o � 7       �����&        �     ��! ���       ���� � ������������}         ����
   " #           L s � :       �����'  �      �     ��! ���       ���� � ������������}         ����
   $ %           P w � =       ����F(  �   	   �     ��! ���       ���� � ������������}         ����
   & '           T { � @       �����(  �      �     ��! ���       ���� � ������������}         ����
   ( )           X  � C       �����)  �#      �	     ��! ���       ���� � ������������}         ����
               D j � .       ����~,  �c      �      ��! ���        ���� � �����  �  ~         ����
               H o � 2       ����P-  �j      �     ��! ���        ���� � �����  �  ~         ����
               L t � 6       ����".  q      �     ��! ���        ���� � �����  �  ~         ����
                P y � :       �����.  �w      �     ��! ���       ���� � �����  �  ~         ����
   ! "           T ~ � >       �����/  0~      �     ��! ���       ���� � �����  �  ~         ����
   $ %           X � � B       �����0  ��   	   �     ��! ���       ���� � �����  �  ~         ����
   & '           \ � � F       ����j1  P�      �     ��! ���       ���� � �����  �  ~         ����
   ( )           ` � J       ����<2  ��      �     ��! ���       ���� � �����  �  ~         ����
   * +           d � 
N       ����3  p�      �     ��! ���       ���� � �����  �  ~         ����
   , -           h � R       �����3   �      �	     ��! ���       ���� � �����  �  ~         ����
               T � � >       ����(7  h�      �      ��! ���        ���� � �����  �           ����
                X � B       ����8  ��      �     ��! ���        ���� � �����  �           ����
   ! "           \ � F       ����9  H      �     ��! ���        ���� � �����  �           ����
   # $           ` � J       �����9  �	   	   �     ��! ���       ���� � �����  �           ����
   % &           d � N       �����:  (      �     ��! ���       ���� � �����  �           ����
   ' (           h � R       �����;  �      �     ��! ���       ���� � �����  �           ����
   * +           l � $V       �����<  #      �     ��! ���       ���� � �����  �           ����
   , -           p � +Z       �����=  x+      �     ��! ���       ���� � �����  �           ����
   . /           t � 2^       �����>  �3      �     ��! ���       ���� � �����  �           ����
   0 1           x � 9b       �����?  X<      �	     ��! ���       ���� � �����  �           ����
   ! "           c � #M       ����XC  p�      �      ��! ���        ����	 � �����  �  �         ����
   # $           g � *Q       ����fD  ��   
   �     ��! ���        ����	 � �����  �  �         ����
   % &           k � 1U       ����tE  ��      �     ��! ���        ����	 � �����  �  �         ����
   ' (           o � 8Y       �����F  �      �     ��! ���       ����	 � �����  �  �         ����
   ) *           s � ?]       �����G  ��      �     ��! ���       ����	 � �����  �  �         ����
   + ,           w � Fa       �����H  ,�      �     ��! ���       ����	 � �����  �  �         ����
   . /           { � Me       �����I  ��      �     ��! ���       ����	 � �����  �  �         ����
   0 1            � Ti       �����J  D�      �     ��! ���       ����	 � �����  �  �         ����
   2 3           � � [m       �����K  ��       �     ��! ���       ����	 � �����  �  �         ����
   4 5           � � bq       �����L  \    ��  �	     ��! ���       ����	 � �����  �  �         ����
   % &           r � K\       ����Q  �{   	   �      ��! ���        ����
 � �����  �  �         ����
   ' (           w � R`       ����:R  ~�      �     ��! ���        ����
 � �����  �  �         ����
   ) *           | � Yd       ����fS  b�      �     ��! ���        ����
 � �����  �  �         ����
   + ,           � � `h       �����T  F�      �     ��! ���       ����
 � �����  �  �         ����
   - .           � � gl       �����U  *�      �     ��! ���       ����
 � �����  �  �         ����
   / 0           � � np       �����V  �      �     ��! ���       ����
 � �����  �  �         ����
   2 3           � � ut       ����X  ��      �     ��! ���       ����
 � �����  �  �         ����
   4 5           � � |x       ����BY  ��   ��  �     ��! ���       ����
 � �����  �  �         ����
   6 7           � � �|       ����nZ  ��   ��  �     ��! ���       ����
 � �����  �  �         ����
   8 9           � � ��       �����[  ��   ��  �	     ��! ���       ����
 �����  �  �         ����
   ) *           � � rj d     ����J`  x�      �      ��! ���        ���� � �����  �  �         ����
   + ,           � � yo e     �����a  �      �     ��! ���        ���� � �����  �  �         ����
   - .           � � �t f     �����b  h�      �     ��! ���        ���� � �����  �  �         ����
   / 0           � � �y g     ����(d  �      �     ��! ���       ���� � �����  �  �         ����
   1 2           � � �~ h     ����re  X�      �     ��! ���       ���� � �����  �  �         ����
   3 4           � � �� i     �����f  ��   ��  �     ��! ���       ���� � �����  �  �         ����
   6 7           � � �� j     ����h  H�   ��  �     ��! ���       ���� � �����  �  �         ����
   8 9           � � �� k     ����Pi  ��   ��  �     ��! ���       ���� � �����  �  �         ����
   : ;           � � �� l     �����j  8�   ��  �     ��! ���       ���� �����  �  �         ����
   < =           � � �� m     �����k  �   ��  �	     ��! ���       ���� �����  �  �         ����
   - .           � � �� n     ����q  ��      �      ��! ���        ���� � �����  �  �         ����
   / 0           � � �� o     ����tr  ��      �     ��! ���        ���� � �����  �  �         ����
   1 2           � � �� p     �����s  ,�      �     ��! ���        ���� � �����  �  �         ����
   3 4           � � �� q     ����Du  t�   ��  �     ��! ���       ���� � �����  �  �         ����
   5 6           � � �� r     �����v  �   ��  �     ��! ���       ���� � �����  �  �         ����
   7 8           � �� s     ����x     ��  �     ��! ���       ���� � �����  �  �         ����
   : ;           � 	�� t     ����|y  L+   ��  �     ��! ���       ����  �����  �  �         ����
   < =           � �� u     �����z  �=   ��  �     ��! ���       ���� �����  �  �         ����
   > ?           � �� v     ����L|  �O   ��  �     ��! ���       ���� �����  �  �         ����
   @ A           � �� w     �����}  $b   ��  �	     ��! ���       ���� �����  �  �         ����
   1 2           � �� x     ����T�  �.      �      ��! ���        ���� � �����  �  �         ����
   3 4           � 	�� y     ����ڄ  �C       �     ��! ���        ���� � �����  �  �         ����
   5 6           � �� z     ����`�  @Y   ��  �     ��! ���        ���� � �����  �  �         ����
   7 8           � �� {     �����  �n   ��  �     ��! ���       ���� � �����  �  �         ����
   9 :           � �� |     ����l�  �   ��  �     ��! ���       ����  �����  �  �         ����
   ; <           � !�� }     �����  <�   ��  �     ��! ���       ���� �����  �  �         ����
   > ?           � '�� ~     ����x�  ��   ��  �     ��! ���       ���� �����  �  �         ����
   @ A           � -��      ������  ��   ��  �     ��! ���       ���� �����  �  �         ����
   B C           � 3� �     ������  8�   ��  �     ��! ���       ���� �����  �  �         ����
   D E           � 9� �     ����
�  ��   ��  �	     ��! ���       ���� #�����  �  �          ����                 / /         �����  X       �      ��! ���        ���� � �������������          ����                 / 4         ����  $       �     ��! ���        ���� � �������������          ����                 / 9         ����0  `       �     ��! ���        ���� � �������������          ����    	             / >         ����N  �       �     ��! ���       ���� � �������������          ����   
              / C         ����l  �       �     ��! ���       ���� � �������������          ����                 / H         �����         �     ��! ���       ���� � �������������          ����                 / M         �����  P       �     ��! ���       ���� � �������������          ����                 / R         �����  �       �     ��! ���       ���� � �������������          ����                 / W         �����  �       �     ��! ���       ���� � �������������          ����                 / \         ����         �	     ��! ���       ���� � �������������          ����                 $ J         ����z  n
       �      ��! ���        ���� � �������������          ����    	             ' O         �����  "       �     ��! ���        ���� � �������������          ����   
              * T         �����  �       �     ��! ���        ���� � �������������          ����                 - Y         ����.  �       �     ��! ���       ���� � �������������          ����                 0 ^         ����j  >       �     ��! ���       ���� � �������������          ����                 3 c         �����  �       �     ��! ���       ���� � �������������          ����                 6 h         �����  �       �     ��! ���       ���� � �������������          ����                 9 m         ����  Z       �     ��! ���       ���� � �������������          ����                 < r         ����Z         �     ��! ���       ���� � �������������          ����                 ? w         �����  �       �	     ��! ���       ���� � �������������         ����   
             + d         �����         �      ��! ���        ���� � �������������         ����               ! / i         �����  �       �     ��! ���        ���� � �������������         ����               $ 3 n         ����:  �       �     ��! ���        ���� � �������������         ����               ' 7 s         �����  P       �     ��! ���       ���� � �������������         ����               * ; x         �����  �       �     ��! ���       ���� � �������������         ����               - ? }         ����H   !       �     ��! ���       ���� � �������������         ����               0 C �         �����  �"       �     ��! ���       ���� � �������������         ����               3 G �         �����  �#       �     ��! ���       ���� � �������������         ����               6 K �         ����V	  X%       �     ��! ���       ���� � �������������         ����               9 O �         �����	  �&       �	     ��! ���       ���� � �������������         ����               & < }        ����  x7       �      ��! ���        ���� � �������������         ����               ) @ �        �����  �9       �     ��! ���        ���� � �������������         ����               , D �         ����  (<       �     ��! ���        ���� � �������������         ����               / H � #       �����  �>       �     ��! ���       ���� � �������������         ����               2 L � &       �����  �@       �     ��! ���       ���� � �������������         ����               5 P � )       ����p  0C       �     ��! ���       ���� � �������������         ����               8 T � ,       �����  �E       �     ��! ���       ���� � �������������         ����               ; X � /       ����`  �G       �     ��! ���       ���� � �������������         ����                > \ � 2       �����  8J       �     ��! ���       ���� � �������������         ����   ! "           A ` � 5       ����P  �L       �	     ��! ���       ���� � �������������         ����               - L � !       ����0   g       �      ��! ���        ���� � �������������         ����               0 P � $       �����  �j       �     ��! ���        ���� � �������������         ����               3 T � '       ����\  (n       �     ��! ���        ���� � �������������         ����               6 X � *       �����  �q       �     ��! ���       ���� � �������������         ����               9 \ � -       �����  0u       �     ��! ���       ���� � �������������         ����               < ` � 0       ����  �x       �     ��! ���       ���� � �������������         ����                ? d � 3       �����  8|       �     ��! ���       ���� � �������������         ����   ! "           B h � 6       ����J  �       �     ��! ���       ���� � �������������         ����   # $           E l � 9       �����  @�    
   �     ��! ���       ���� � �������������         ����   % &           H p � <       ����v  Ć    	   �	     ��! ���       ���� � �������������         ����               4 [ � (       �����  ��       �      ��! ���        ���� � �������������         ����               8 _ � +       �����  ��       �     ��! ���        ���� � �������������         ����               < c � .       ����6  z�       �     ��! ���        ���� � �������������         ����               @ g � 1       �����  f�       �     ��! ���       ���� � �������������         ����               D k � 4       �����  R�       �     ��! ���       ���� � �������������         ����   ! "           H o � 7       ����R  >�       �     ��! ���       ���� � �������������         ����   # $           L s � :       ����  *�       �     ��! ���       ���� � �������������         ����   % &           P w � =       �����  �    	   �     ��! ���       ���� � �������������         ����   ' (           T { � @       ����n  �       �     ��! ���       ���� � �������������         ����   ) *           X  � C       ����"  ��       �	     ��! ���       ���� � �������������         ����               D j � .       �����!  �      �      ��! ���        ���� � �����  �  �         ����               H o � 2       �����"         �     ��! ���        ���� � �����  �  �         ����               L t � 6       �����#  �      �     ��! ���        ���� � �����  �  �         ����     !           P y � :       ����h$  @#      �     ��! ���       ���� � �����  �  �         ����   " #           T ~ � >       ����:%  �)      �     ��! ���       ���� � �����  �  �         ����   $ %           X �  B       ����&  `0   	   �     ��! ���       ���� � �����  �  �         ����   ' (           \ � F       �����&  �6      �     ��! ���       ���� � �����  �  �         ����   ) *           ` � J       �����'  �=      �     ��! ���       ���� � �����  �  �         ����   + ,           d � N       �����(  D      �     ��! ���       ���� � �����  �  �         ����   - .           h � R       ����T)  �J      �	     ��! ���       ���� � �����  �  �         ����               T � >       �����,  |�      �      ��! ���        ���� � �����  �  �         ����     !           X � 	B       �����-  �      �     ��! ���        ���� � �����  �  �         ����   " #           \ � F       ����|.  \�      �     ��! ���        ���� � �����  �  �         ����   $ %           ` � J       ����l/  ̪   	   �     ��! ���       ���� � �����  �  �         ����   & '           d � N       ����\0  <�      �     ��! ���       ���� � �����  �  �         ����   ( )           h � %R       ����L1  ��      �     ��! ���       ���� � �����  �  �         ����   + ,           l � ,V       ����<2  �      �     ��! ���       ���� � �����  �  �         ����   - .           p � 3Z       ����,3  ��      �     ��! ���       ���� � �����  �  �         ����   / 0           t � :^       ����4  ��      �     ��! ���       ���� � �����  �  �         ����   1 2           x � Ab       ����5  l�      �	     ��! ���       ���� � �����  �  �         ����   " #           c � +M       �����8  �7      �      ��! ���        ����	 � �����  �  �         ����   $ %           g � 2Q       �����9  �B   
   �     ��! ���        ����	 � �����  �  �         ����   & '           k � 9U       �����:  M      �     ��! ���        ����	 � �����  �  �         ����   ( )           o � @Y       �����;  �W      �     ��! ���       ����	 � �����  �  �         ����   * +           s � G]       ����=  (b      �     ��! ���       ����	 � �����  �  �         ����   , -           w � Na       ����>  �l      �     ��! ���       ����	 � �����  �  �         ����   / 0           { � Ue       ���� ?  @w      �     ��! ���       ����	 � �����  �  �         ����   1 2            � \i       ����.@  ́      �     ��! ���       ����	 � �����  �  �         ����   3 4           � � cm       ����<A  X�       �     ��! ���       ����	 � �����  �  �         ����   5 6           � � jq       ����JB  �   ��  �	     ��! ���       ����	 � �����  �  �         ����   & '           r � S\       �����F  �   	   �      ��! ���        ����
 � �����  �  �         ����   ( )           w � Z`       �����G  z      �     ��! ���        ����
 � �����  �  �         ����   * +           | � ad       �����H  ^!      �     ��! ���        ����
 � �����  �  �         ����   , -           � � hh       ����J  B.      �     ��! ���       ����
 � �����  �  �         ����   . /           � � ol       ����2K  &;      �     ��! ���       ����
 � �����  �  �         ����   0 1           � � vp       ����^L  
H      �     ��! ���       ����
 � �����  �  �         ����   3 4           � � }t       �����M  �T      �     ��! ���       ����
 � �����  �  �         ����   5 6           � � �x       �����N  �a   ��  �     ��! ���       ����
 � �����  �  �         ����   7 8           � � �|       �����O  �n   ��  �     ��! ���       ����
 � �����  �  �         ����   9 :           � � ��       ����Q  �{   ��  �	     ��! ���       ����
 �����  �  �         ����   * +           � � zj d     �����U  �      �      ��! ���        ���� � �����  �  �         ����   , -           � � �o e     ����W  `      �     ��! ���        ���� � �����  �  �         ����   . /           � � �t f     ����RX  �#      �     ��! ���        ���� � �����  �  �         ����   0 1           � � �y g     �����Y  P3      �     ��! ���       ���� � �����  �  �         ����   2 3           � � �~ h     �����Z  �B      �     ��! ���       ���� � �����  �  �         ����   4 5           � � �� i     ����0\  @R   ��  �     ��! ���       ���� � �����  �  �         ����   7 8           � � �� j     ����z]  �a   ��  �     ��! ���       ���� � �����  �  �         ����   9 :           � � �� k     �����^  0q   ��  �     ��! ���       ���� � �����  �  �         ����   ; <           � � �� l     ����`  ��   ��  �     ��! ���       ���� �����  �  �         ����   = >           � � �� m     ����Xa   �   ��  �	     ��! ���       ���� �����  �  �         ����   . /           � � �� n     �����f  �4      �      ��! ���        ���� � �����  �  �         ����   0 1           � � �� o     �����g  �F      �     ��! ���        ���� � �����  �  �         ����   2 3           � � �� p     ����Pi  Y      �     ��! ���        ���� � �����  �  �         ����   4 5           � � �� q     �����j  Xk   ��  �     ��! ���       ���� � �����  �  �         ����   6 7           � � �� r     ���� l  �}   ��  �     ��! ���       ���� � �����  �  �         ����   8 9           � �� s     �����m  �   ��  �     ��! ���       ���� � �����  �  �         ����   ; <           � 	�� t     �����n  0�   ��  �     ��! ���       ����  �����  �  �         ����   = >           � �� u     ����Xp  x�   ��  �     ��! ���       ���� �����  �  �         ����   ? @           � �� v     �����q  ��   ��  �     ��! ���       ���� �����  �  �         ����   A B           � �� w     ����(s  �   ��  �	     ��! ���       ���� �����  �  �         ����   2 3           � �� x     �����x  �      �      ��! ���        ���� � �����  �  �         ����   4 5           � 	�� y     ����Nz  D�       �     ��! ���        ���� � �����  �  �         ����   6 7           � �� z     �����{  ��   ��  �     ��! ���        ���� � �����  �  �         ����   8 9           � �� {     ����Z}  ��   ��  �     ��! ���       ���� � �����  �  �         ����   : ;           � �� |     �����~  @�   ��  �     ��! ���       ����  �����  �  �         ����   < =           � !�� }     ����f�  �   ��  �     ��! ���       ���� �����  �  �         ����   ? @           � '�� ~     �����  �   ��  �     ��! ���       ���� �����  �  �         ����   A B           � -�      ����r�  <0   ��  �     ��! ���       ���� �����  �  �         ����   C D           � 3� �     ������  �E   ��  �     ��! ���       ���� �����  �  �         ����   E F           � 9� �     ����~�  �Z   ��  �	     ��! ���       ���� #�����  �  �          ����                 7 7         �����  �        6      ��! ���        ���� � �������������          ����                 7 <         �����  |       6     ��! ���        ���� � �������������          ����                 7 A         �����  �       6     ��! ���        ���� � �������������          ����    	             7 F         �����  �       6     ��! ���       ���� � �������������          ����   
              7 K         ����  0        6     ��! ���       ���� � �������������          ����                 7 P         ����6  l        6     ��! ���       ���� � �������������          ����                 7 U         ����T  �        6     ��! ���       ���� � �������������          ����                 7 Z         ����r  �        6     ��! ���       ���� � �������������          ����                 7 _         �����   !       6     ��! ���       ���� � �������������          ����                 7 d         �����  \!       6	     ��! ���       ���� � �������������          ����                 $ R         ����&  r3       7      ��! ���        ���� � �������������          ����    	             ' W         ����b  &4       7     ��! ���        ���� � �������������          ����   
              * \         �����  �4       7     ��! ���        ���� � �������������          ����                 - a         �����  �5       7     ��! ���       ���� � �������������          ����                 0 f         ����  B6       7     ��! ���       ���� � �������������          ����                 3 k         ����R  �6       7     ��! ���       ���� � �������������          ����                 6 p         �����  �7       7     ��! ���       ���� � �������������          ����                 9 u         �����  ^8       7     ��! ���       ���� � �������������          ����                 < z         ����  9       7     ��! ���       ���� � �������������          ����                 ?          ����B  �9       7	     ��! ���       ���� � �������������         ����   
             + l         ����2  �P       8      ��! ���        ���� � �������������         ����               ! / q         �����  0R       8     ��! ���        ���� � �������������         ����               $ 3 v         �����  �S       8     ��! ���        ���� � �������������         ����               ' 7 {         ����@   U       8     ��! ���       ���� � �������������         ����               * ; �         �����  hV       8     ��! ���       ���� � �������������         ����               - ? �         �����  �W       8     ��! ���       ���� � �������������         ����               0 C �         ����N  8Y       8     ��! ���       ���� � �������������         ����               3 G �         �����  �Z       8     ��! ���       ���� � �������������         ����               6 K �         ����  \       8     ��! ���       ���� � �������������         ����               9 O �         ����\  p]       8	     ��! ���       ���� � �������������         ����               & < �        �����  �{       9      ��! ���        ���� � �������������         ����               ) @ �        ����<  ,~       9     ��! ���        ���� � �������������         ����               , D �         �����  ��       9     ��! ���        ���� � �������������         ����               / H � #       ����,  ܂       9     ��! ���       ���� � �������������         ����               2 L � &       �����  4�       9     ��! ���       ���� � �������������         ����               5 P � )       ����  ��       9     ��! ���       ���� � �������������         ����               8 T � ,       �����  �       9     ��! ���       ���� � �������������         ����               ; X � /       ����  <�       9     ��! ���       ���� � �������������         ����                > \ � 2       �����  ��       9     ��! ���       ���� � �������������         ����   ! "           A ` � 5       �����  �       9	     ��! ���       ���� � �������������         ����               - L � !       �����  (�       :      ��! ���        ���� � �������������         ����               0 P � $       ����r  ��       :     ��! ���        ���� � �������������         ����               3 T � '       ����   0�       :     ��! ���        ���� � �������������         ����               6 X � *       �����   ��       :     ��! ���       ���� � �������������         ����               9 \ � -       ����4!  8�       :     ��! ���       ���� � �������������         ����               < ` � 0       �����!  ��       :     ��! ���       ���� � �������������         ����                ? d � 3       ����`"  @�       :     ��! ���       ���� � �������������         ����   ! "           B h � 6       �����"  ��       :     ��! ���       ���� � �������������         ����   # $           E l � 9       �����#  H�    
   :     ��! ���       ���� � �������������         ����   % &           H p � <       ����"$  ��    	   :	     ��! ���       ���� � �������������         ����               4 [ � (       ����z&  V      ;      ��! ���        ���� � �������������         ����               8 _ � +       ����.'  B      ;     ��! ���        ���� � �������������         ����               < c � .       �����'  .      ;     ��! ���        ���� � �������������         ����               @ g � 1       �����(        ;     ��! ���       ���� � �������������         ����               D k � 4       ����J)  !      ;     ��! ���       ���� � �������������         ����   ! "           H o � 7       �����)  �%      ;     ��! ���       ���� � �������������         ����   # $           L s � :       �����*  �*      ;     ��! ���       ���� � �������������         ����   % &           P w � =       ����f+  �/   	   ;     ��! ���       ���� � �������������         ����   ' (           T { � @       ����,  �4      ;     ��! ���       ���� � �������������         ����   ) *           X  � C       �����,  �9      ;	     ��! ���       ���� � �������������         ����               D j � .       �����/  �|      <      ��! ���        ���� � �����  �  �         ����               H o � 2       ����p0  ��      <     ��! ���        ���� � �����  �  �         ����               L t � 6       ����B1  �      <     ��! ���        ���� � �����  �  �         ����     !           P y � :       ����2  ��      <     ��! ���       ���� � �����  �  �         ����   " #           T ~ >       �����2  0�      <     ��! ���       ���� � �����  �  �         ����   $ %           X � B       �����3  ��   	   <     ��! ���       ���� � �����  �  �         ����   ' (           \ � F       �����4  P�      <     ��! ���       ���� � �����  �  �         ����   ) *           ` � J       ����\5  �      <     ��! ���       ���� � �����  �  �         ����   + ,           d � N       ����.6  p�      <     ��! ���       ���� � �����  �  �         ����   - .           h �  R       ���� 7   �      <	     ��! ���       ���� � �����  �  �         ����               T � 
>       ����H:  �      =      ��! ���        ���� � �����  �  �         ����     !           X � B       ����8;  �      =     ��! ���        ���� � �����  �  �         ����   " #           \ � F       ����(<  h      =     ��! ���        ���� � �����  �  �         ����   $ %           ` � J       ����=  �%   	   =     ��! ���       ���� � �����  �  �         ����   & '           d � &N       ����>  H.      =     ��! ���       ���� � �����  �  �         ����   ( )           h � -R       �����>  �6      =     ��! ���       ���� � �����  �  �         ����   + ,           l � 4V       �����?  (?      =     ��! ���       ���� � �����  �  �         ����   - .           p � ;Z       �����@  �G      =     ��! ���       ���� � �����  �  �         ����   / 0           t � B^       �����A  P      =     ��! ���       ���� � �����  �  �         ����   1 2           x � Ib       �����B  xX      =	     ��! ���       ���� � �����  �  �         ����   " #           c � 3M       ����xF  ��      >      ��! ���        ����	 � �����  �  �         ����   $ %           g � :Q       �����G  <�   
   >     ��! ���        ����	 � �����  �  �         ����   & '           k � AU       �����H  ��      >     ��! ���        ����	 � �����  �  �         ����   ( )           o � HY       �����I  T�      >     ��! ���       ����	 � �����  �  �         ����   * +           s � O]       �����J  ��      >     ��! ���       ����	 � �����  �  �         ����   , -           w � Va       �����K  l�      >     ��! ���       ����	 � �����  �  �         ����   / 0           { � ]e       �����L  ��      >     ��! ���       ����	 � �����  �  �         ����   1 2            � di       �����M  �
      >     ��! ���       ����	 � �����  �  �         ����   3 4           � � km       �����N         >     ��! ���       ����	 � �����  �  �         ����   5 6           � � rq       �����O  �   ��  >	     ��! ���       ����	 � �����  �  �         ����   & '           r � [\       ����.T  ��   	   ?      ��! ���        ����
 � �����  �  �         ����   ( )           w � b`       ����ZU  ު      ?     ��! ���        ����
 � �����  �  �         ����   * +           | � id       �����V  ·      ?     ��! ���        ����
 � �����  �  �         ����   , -           � � ph       �����W  ��      ?     ��! ���       ����
 � �����  �  �         ����   . /           � � wl       �����X  ��      ?     ��! ���       ����
 � �����  �  �         ����   0 1           � � ~p       ����
Z  n�      ?     ��! ���       ����
 � �����  �  �         ����   3 4           � � �t       ����6[  R�      ?     ��! ���       ����
 � �����  �  �         ����   5 6           � � �x       ����b\  6�   ��  ?     ��! ���       ����
 � �����  �  �         ����   7 8           � � �|       �����]     ��  ?     ��! ���       ����
 � �����  �  �         ����   9 :           � � ��       �����^  �   ��  ?	     ��! ���       ����
 �����  �  �         ����   * +           � � �j d     ����jc  ��      @      ��! ���        ���� � �����  �  �         ����   , -           � � �o e     �����d  p�      @     ��! ���        ���� � �����  �  �         ����   . /           � � �t f     �����e  ��      @     ��! ���        ���� � �����  �  �         ����   0 1           � � �y g     ����Hg  `�      @     ��! ���       ���� � �����  �  �         ����   2 3           � � �~ h     �����h  ��      @     ��! ���       ���� � �����  �  �         ����   4 5           � � �� i     �����i  P�   ��  @     ��! ���       ���� � �����  �  �         ����   7 8           � � �� j     ����&k  �   ��  @     ��! ���       ���� � �����  �  �         ����   9 :           � � �� k     ����pl  @   ��  @     ��! ���       ���� � �����  �  �         ����   ; <           � � �� l     �����m  �$   ��  @     ��! ���       ���� �����  �  �         ����   = >           � � �� m     ����o  04   ��  @	     ��! ���       ���� �����  �  �         ����   . /           � � �� n     ����,t  <�      A      ��! ���        ���� � �����  �  �         ����   0 1           � � �� o     �����u  ��      A     ��! ���        ���� � �����  �  �         ����   2 3           � � �� p     �����v  �
      A     ��! ���        ���� � �����  �  �         ����   4 5           � � �� q     ����dx     ��  A     ��! ���       ���� � �����  �  �         ����   6 7           � � �� r     �����y  \/   ��  A     ��! ���       ���� � �����  �  �         ����   8 9           � �� s     ����4{  �A   ��  A     ��! ���       ���� � �����  �  �         ����   ; <           � 	�� t     �����|  �S   ��  A     ��! ���       ����  �����  �  �         ����   = >           � �� u     ����~  4f   ��  A     ��! ���       ���� �����  �  �         ����   ? @           � �� v     ����l  |x   ��  A     ��! ���       ���� �����  �  �         ����   A B           � �� w     ����Ԁ  Ċ   ��  A	     ��! ���       ���� �����  �  �         ����   2 3           � �� x     ����t�  XZ      B      ��! ���        ���� � �����  �  �         ����   4 5           � 	�� y     ������  �o       B     ��! ���        ���� � �����  �  �         ����   6 7           � �� z     ������   �   ��  B     ��! ���        ���� � �����  �  �         ����   8 9           � �� {     �����  T�   ��  B     ��! ���       ���� � �����  �  �         ����   : ;           � �� |     ������  ��   ��  B     ��! ���       ����  �����  �  �         ����   < =           � !�� }     �����  ��   ��  B     ��! ���       ���� �����  �  �         ����   ? @           � '� ~     ������  P�   ��  B     ��! ���       ���� �����  �  �         ����   A B           � -�      �����  ��   ��  B     ��! ���       ���� �����  �  �         ����   C D           � 3� �     ������  �   ��  B     ��! ���       ���� �����  �  �         ����   E F           � 9� �     ����*�  L   ��  B	     ��! ���       ���� #�����  �  �          ����                 9 9         ����0  �        �      ��! ���        ���� � �������������          ����                 9 >         ����N  �"       �     ��! ���        ���� � �������������          ����                 9 C         ����l  �"       �     ��! ���        ���� � �������������          ����    	             9 H         �����  #       �     ��! ���       ���� � �������������          ����   
              9 M         �����  P#       �     ��! ���       ���� � �������������          ����                 9 R         �����  �#       �     ��! ���       ���� � �������������          ����                 9 W         �����  �#       �     ��! ���       ���� � �������������          ����                 9 \         ����  $       �     ��! ���       ���� � �������������          ����                 9 a         ����   @$       �     ��! ���       ���� � �������������          ����                 9 f         ����>  |$       �	     ��! ���       ���� � �������������          ����                 $ V         �����  "8       �      ��! ���        ���� � �������������          ����    	             ' [         �����  �8       �     ��! ���        ���� � �������������          ����   
              * `         ����.  �9       �     ��! ���        ���� � �������������          ����                 - e         ����j  >:       �     ��! ���       ���� � �������������          ����                 0 j         �����  �:       �     ��! ���       ���� � �������������          ����                 3 o         �����  �;       �     ��! ���       ���� � �������������          ����                 6 t         ����  Z<       �     ��! ���       ���� � �������������          ����                 9 y         ����Z  =       �     ��! ���       ���� � �������������          ����                 < ~         �����  �=       �     ��! ���       ���� � �������������          ����                 ? �         �����  v>       �	     ��! ���       ���� � �������������         ����   
             + r         �����  W       �      ��! ���        ���� � �������������         ����               ! / w         ����  pX       �     ��! ���        ���� � �������������         ����               $ 3 |         ����v  �Y       �     ��! ���        ���� � �������������         ����               ' 7 �         �����  @[       �     ��! ���       ���� � �������������         ����               * ; �         ����*  �\       �     ��! ���       ���� � �������������         ����               - ? �         �����  ^       �     ��! ���       ���� � �������������         ����               0 C �         �����  x_       �     ��! ���       ���� � �������������         ����               3 G �         ����8  �`       �     ��! ���       ���� � �������������         ����               6 K �         �����  Hb       �     ��! ���       ���� � �������������         ����               9 O �         �����  �c       �	     ��! ���       ���� � �������������         ����               # ; �        ����T  ��       �      ��! ���        ���� � �������������         ����               & ? �        �����  ��       �     ��! ���        ���� � �������������         ����               ) C �         ����D  T�       �     ��! ���        ���� � �������������         ����               , G � #       �����  ��       �     ��! ���       ���� � �������������         ����               / K � &       ����4  �       �     ��! ���       ���� � �������������         ����               2 O � )       �����  \�       �     ��! ���       ���� � �������������         ����               5 S � ,       ����$  ��       �     ��! ���       ���� � �������������         ����               8 W � /       �����  �       �     ��! ���       ���� � �������������         ����                ; [ � 2       ����  d�       �     ��! ���       ���� � �������������         ����   ! "           > _ � 5       �����  ��       �	     ��! ���       ���� � �������������         ����               ' J � !       ����l   ��       �      ��! ���        ���� � �������������         ����               * N � $       ����!  �       �     ��! ���        ���� � �������������         ����               - R � '       �����!  ��       �     ��! ���        ���� � �������������         ����               0 V � *       ����."  �       �     ��! ���       ���� � �������������         ����               3 Z � -       �����"  ��       �     ��! ���       ���� � �������������         ����               6 ^ � 0       ����Z#  �       �     ��! ���       ���� � �������������         ����                9 b � 3       �����#  ��       �     ��! ���       ���� � �������������         ����   ! "           < f � 6       �����$  $�       �     ��! ���       ���� � �������������         ����   # $           ? j � 9       ����%  ��    
   �     ��! ���       ���� � �������������         ����   % &           B n � <       �����%  ,�    	   �	     ��! ���       ���� � �������������         ����               + Y � (       ����
(  F      �      ��! ���        ���� � �������������         ����               / ] � +       �����(  2      �     ��! ���        ���� � �������������         ����               3 a � .       ����r)  "      �     ��! ���        ���� � �������������         ����               7 e � 1       ����&*  
'      �     ��! ���       ���� � �������������         ����               ; i � 4       �����*  �+      �     ��! ���       ���� � �������������         ����   ! "           ? m � 7       �����+  �0      �     ��! ���       ���� � �������������         ����   # $           C q � :       ����B,  �5      �     ��! ���       ���� � �������������         ����   % &           G u =       �����,  �:   	   �     ��! ���       ���� � �������������         ����   ' (           K y @       �����-  �?      �     ��! ���       ���� � �������������         ����   ) *           O } C       ����^.  �D      �	     ��! ���       ���� � �������������         ����               8 g � .       ����.1  p�      �      ��! ���        ���� � �����  �  �         ����               < l 2       ���� 2   �      �     ��! ���        ���� � �����  �  �         ����               @ q 6       �����2  ��      �     ��! ���        ���� � �����  �  �         ����     !           D v :       �����3   �      �     ��! ���       ���� � �����  �  �         ����   " #           H { >       ����v4  ��      �     ��! ���       ���� � �����  �  �         ����   $ %           L � B       ����H5  @�   	   �     ��! ���       ���� � �����  �  �         ����   ' (           P �  F       ����6  а      �     ��! ���       ���� � �����  �  �         ����   ) *           T � &J       �����6  `�      �     ��! ���       ���� � �����  �  �         ����   + ,           X � ,N       �����7  �      �     ��! ���       ���� � �����  �  �         ����   - .           \ � 2R       �����8  ��      �	     ��! ���       ���� � �����  �  �         ����               D ~  >       �����;  �      �      ��! ���        ���� � �����  �  �         ����     !           H � 'B       �����<  #      �     ��! ���        ���� � �����  �  �         ����   " #           L � .F       �����=  x+      �     ��! ���        ���� � �����  �  �         ����   $ %           P � 5J       �����>  �3   	   �     ��! ���       ���� � �����  �  �         ����   & '           T � <N       �����?  X<      �     ��! ���       ���� � �����  �  �         ����   ( )           X � CR       �����@  �D      �     ��! ���       ���� � �����  �  �         ����   + ,           \ � JV       ����xA  8M      �     ��! ���       ���� � �����  �  �         ����   - .           ` � QZ       ����hB  �U      �     ��! ���       ���� � �����  �  �         ����   / 0           d � X^       ����XC  ^      �     ��! ���       ���� � �����  �  �         ����   1 2           h � _b       ����HD  �f      �	     ��! ���       ���� � �����  �  �         ����   " #           O � MM       ����H  P�      �      ��! ���        ����	 � �����  �  �         ����   $ %           S � TQ       ����I  ��   
   �     ��! ���        ����	 � �����  �  �         ����   & '           W � [U       ����$J  h�      �     ��! ���        ����	 � �����  �  �         ����   ( )           [ � bY       ����2K  ��      �     ��! ���       ����	 � �����  �  �         ����   * +           _ � i]       ����@L  ��      �     ��! ���       ����	 � �����  �  �         ����   , -           c � pa       ����NM        �     ��! ���       ����	 � �����  �  �         ����   / 0           g � we       ����\N  �      �     ��! ���       ����	 � �����  �  �         ����   1 2           k � ~i       ����jO  $      �     ��! ���       ����	 � �����  �  �         ����   3 4           o � �m       ����xP  �$       �     ��! ���       ����	 � �����  �  �         ����   5 6           s � �q       �����Q  </   ��  �	     ��! ���       ����	 � �����  �  �         ����   & '           Y � z\       �����U  *�   	   �      ��! ���        ����
 � �����  �  �         ����   ( )           ^ � �`       �����V  �      �     ��! ���        ����
 � �����  �  �         ����   * +           c � �d       ����X  ��      �     ��! ���        ����
 � �����  �  �         ����   , -           h � �h       ����BY  ��      �     ��! ���       ����
 � �����  �  �         ����   . /           m � �l       ����nZ  ��      �     ��! ���       ����
 � �����  �  �         ����   0 1           r � �p       �����[  ��      �     ��! ���       ����
 � �����  �  �         ����   3 4           w � �t       �����\  ��      �     ��! ���       ����
 � �����  �  �         ����   5 6           | � �x       �����]  f	   ��  �     ��! ���       ����
 � �����  �  �         ����   7 8           � � �|       ����_  J   ��  �     ��! ���       ����
 � �����  �  �         ����   9 :           � � ��       ����J`  .#   ��  �	     ��! ���       ����
 �����  �  �         ����   * +           l � �j d     �����d  ��      �      ��! ���        ���� � �����  �  �         ����   , -           q � �o e     ����Df  0�      �     ��! ���        ���� � �����  �  �         ����   . /           v � �t f     �����g  ��      �     ��! ���        ���� � �����  �  �         ����   0 1           { � �y g     �����h   �      �     ��! ���       ���� � �����  �  �         ����   2 3           � � �~ h     ����"j  ��      �     ��! ���       ���� � �����  �  �         ����   4 5           � � �� i     ����lk  	   ��  �     ��! ���       ���� � �����  �  �         ����   7 8           � � �� j     �����l  �   ��  �     ��! ���       ���� � �����  �  �         ����   9 :           � � �� k     ���� n   (   ��  �     ��! ���       ���� � �����  �  �         ����   ; <           � � �� l     ����Jo  x7   ��  �     ��! ���       ���� �����  �  �         ����   = >           � � �� m     �����p  �F   ��  �	     ��! ���       ���� �����  �  �         ����   . /           ~ � �� n     �����u  ��      �      ��! ���        ���� � �����  �  �         ����   0 1           � � �� o     ����$w  �      �     ��! ���        ���� � �����  �  �         ����   2 3           � � �� p     �����x        �     ��! ���        ���� � �����  �  �         ����   4 5           � � �� q     �����y  d1   ��  �     ��! ���       ���� � �����  �  �         ����   6 7           � � �� r     ����\{  �C   ��  �     ��! ���       ���� � �����  �  �         ����   8 9           � � �� s     �����|  �U   ��  �     ��! ���       ���� � �����  �  �         ����   ; <           � � t     ����,~  <h   ��  �     ��! ���       ����  �����  �  �         ����   = >           � 
� u     �����  �z   ��  �     ��! ���       ���� �����  �  �         ����   ? @           � � v     ������  ̌   ��  �     ��! ���       ���� �����  �  �         ����   A B           � � w     ����d�  �   ��  �	     ��! ���       ���� �����  �  �         ����   2 3           � � � x     �����  8p      �      ��! ���        ���� � �����  �  �         ����   4 5           �  � y     ������  ��       �     ��! ���        ���� � �����  �  �         ����   6 7           � � z     �����  ��   ��  �     ��! ���        ���� � �����  �  �         ����   8 9           � � {     ������  4�   ��  �     ��! ���       ���� � �����  �  �         ����   : ;           � '� |     �����  ��   ��  �     ��! ���       ����  �����  �  �         ����   < =           � /� }     ������  ��   ��  �     ��! ���       ���� �����  �  �         ����   ? @           � 7� ~     ����(�  0�   ��  �     ��! ���       ���� �����  �  �         ����   A B           � $?�      ������  �   ��  �     ��! ���       ���� �����  �  �         ����   C D           � *G� �     ����4�  �   ��  �     ��! ���       ���� �����  �  �         ����   E F           � 0O� �     ������  ,0   ��  �	     ��! ���       ���� #�����  �  �         ����    1 2            � �         	      �        �        ��         ����c   �������������         ����    3 4            � �            >  |        �       ��         ����c   �������������         ����    5 6            � �            \  �        �       ��         ����c   �������������         ����    7 8            � �            z  �        �       ��        ����c   �������������         ����    9 :            � �            �  0        �       ��        ����c   �������������         ����    ; <            � �            �  l        �       ��        ����c   �������������         ����    = >            � �            �  �        �       ��        ����c   �������������         ����    ? @            � �            �  �        �       ��        ����c   �������������         ����    A B            � �                       �       ��        ����c   �������������         ����    C D            � �            .  \        �	       ��        ����c   �������������         ����   0 1            � �            ,  h        �        ��        ����c   �������������         ����   2 3            � �            J  �        �       ��        ����c   �������������         ����   4 5            � �            h  �        �       ��        ����c   �������������         ����   6 7            � �            �          �       ��       ����c   �������������         ����   8 9            � �            �  H        �       ��       ����c   �������������         ����   : ;            � �         	   �  �        �       ��       ����c   �������������         ����   < =            � �         	   �  �        �       ��       ����c   �������������         ����   > ?            � �         
   �  �        �       ��       ����c   �������������         ����   @ A            � �         
     8        �       ��       ����c   �������������         ����   B C            � �            :  t        �	       ��       ����c   �������������         ����   0 1            � �            �   �         T        ��        ����c   �������������         ����   2 3            � �            �   �        T       ��        ����c   �������������         ����   4 5            � �                      T       ��        ����c   �������������         ����   6 7            � �            "  D        T       ��       ����c   �������������         ����   8 9            � �            @  �        T       ��       ����c   �������������         ����   : ;            � �            ^  �        T       ��       ����c   �������������         ����   < =            � �            |  �        T       ��       ����c   �������������         ����   > ?            � �            �  4        T       ��       ����c   �������������         ����   @ A            � �            �  p        T       ��       ����c   �������������         ����   B C            � �         	   �  �        T	       ��       ����c   �������������         ����   1 2            � �         !   �  /        �        ��        ����c   �������������         ����   3 4            � �         (   �  �        �       ��        ����c   �������������         ����   5 6            � �         )             �       ��        ����c   �������������         ����   7 8            � �         )   *  T        �       ��       ����c   �������������         ����   9 :            � �         *   H  �        �       ��       ����c   �������������         ����   ; <            � �         +   f  �        �       ��       ����c   �������������         ����   = >            � �         +   �          �       ��       ����c   �������������         ����   ? @            � �         ,   �  D        �       ��       ����c   �������������         ����   A B            � �         ,   �  �        �       ��       ����c   �������������         ����   C D            � �         -   �  �        �	       ��       ����c   �������������         ����   1 2            � �            @  �                 ��        ����c   �������������         ����   3 4            � �             ^  �                ��        ����c   �������������         ����   5 6            � �         !   |  �                ��        ����c   �������������         ����   7 8            � �         !   �  4                ��       ����c   �������������         ����   9 :            � �         "   �  p                ��       ����c   �������������         ����   ; <            � �         #   �  �                ��       ����c   �������������         ����   = >            � �         #   �  �                ��       ����c   �������������         ����   ? @            � �         $     $                ��       ����c   �������������         ����   A B            � �         $   0  `                ��       ����c   �������������         ����   C D            � �         %   N  �         	       ��       ����c   �������������         ����   0 1            � �            �  F        �        ��        ����c   �������������         ����   2 3            � �            �  �	        �       ��        ����c   �������������         ����   4 5            � �            �  �	        �       ��        ����c   �������������         ����   6 7            � �            
  
        �       ��       ����c   �������������         ����   8 9            � �            (  P
        �       ��       ����c   �������������         ����   : ;            � �            F  �
        �       ��       ����c   �������������         ����   < =            � �            d  �
        �       ��       ����c   �������������         ����   > ?            � �            �          �       ��       ����c   �������������         ����   @ A            � �            �  @        �       ��       ����c   �������������         ����   B C            � �            �  |        �	       ��       ����c   �������������         ����   1 2            � �         2   `	  �        �      �           ����c   �������������         ����   3 4            � �         0   ~	  �        �     �           ����c   �������������         ����   5 6            � �         1   �	  8        �     �           ����c   �������������         ����   7 8            � �         1   �	  t        �     �          ����c   �������������         ����   9 :            � �         2   �	  �        �     �          ����c   �������������         ����   ; <            � �         3   �	  �        �     �          ����c   �������������         ����   = >            � �         3   
  (        �     �          ����c   �������������         ����   ? @            � �         4   2
  d        �     �          ����c   �������������         ����   A B            � �         4   P
  �        �     �          ����c   �������������         ����   C D            � �         5   n
  �        �	     �          ����c   �������������         ����� ��                            �����  �       L      ��Y ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��	        ������  ����������������       ����� ��                            ����'   N        �      ��R ��
        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������          ���/�/2    ,d d 2           0  �        @       >       �������c   �������������            ���J�J2    1i i 7           N  �        @      >       �������c   �������������            ���e�e2    6n n <           l  �        @      >       �������c   �������������            ������2    ;s s A           �          @      >      �������c   �������������            ������2    @x x F           �  P        @      >      �������c   �������������            ����2    E} } K           �  �        @      >      �������c   �������������            ��)�)�2    J� � P           �  �        @      >      �������c   �������������            ��C�C�2    O� � U                     @      >      �������c   �������������            ��]]2    T� � Z              @        @      >      �������c   �������������            ��w"w"2    Y� � _           >  |        @ 	     >      �������c   �������������            �����2    ,d d 2           �          V       S       �������c   �������������            ��'��2    1i i 7           �  �        V      S       �������c   �������������            ��C�+�2    6n n <           �  �        V      S       �������c   �������������            ��_C�2    ;s s A                     V      S      �������c   �������������            ��{![�2    @x x F              @        V      S      �������c   �������������            ���>s2    E} } K           >  |        V      S      �������c   �������������            ���[�12    J� � P           \  �        V      S      �������c   �������������            ���x�K2    O� � U           z  �        V      S      �������c   �������������            �����e2    T� � Z           �  0        V      S      �������c   �������������            ����2    Y� � _           �  l        V 	     S      �������c   �������������            ���/�T2    d d ,2           �
  L6        o       k       �������c   �������������            ���G�s2    i i 17           T  �8        o      k       �������c   �������������            ���_��2    n n 6<           �  �:        o      k       �������c   �������������            ���w�2    s s ;A           D  T=        o      k      �������c   �������������            ����3�2    x x @F           �  �?        o      k      �������c   �������������            ����Q�2    } } EK           4  B        o      k      �������c   �������������            ���o2    � � JP           �  \D        o      k      �������c   �������������            ��#��-2    � � OU           $  �F        o      k      �������c   �������������            ��:��L2    � � TZ           �  I        o      k      �������c   �������������            ��Q�k2    � � Y_             dK        o 	     k      �������c   �������������             S�S�
2    ,d d 2           �  �        �       �       �������c   �������������             l
l

2    1i i 7           X  `        �      �       �������c   �������������             �%�%
2    6n n <           �  �        �      �       �������c   �������������             �@�@
2    ;s s A             0         �      �      �������c   �������������             �[�[
2    @x x F           f  �!        �      �      �������c   �������������             �v�v
2    E} } K           �   #        �      �      �������c   �������������             ����
2    J� � P           	  h$        �      �      �������c   �������������             ��
2    O� � U           t	  �%        �      �      �������c   �������������             ��
2    T� � Z           �	  8'        �      �      �������c   �������������             4�4�
2    Y� � _           (
  �(        � 	     �      �������c   �������������             a�/2    d ,d 2           j  >        �       �       �������c   �������������             ~6�G2    i 1i 7           �  �        �      �       �������c   �������������             �T�_2    n 6n <           �  �        �      �       �������c   �������������             �r�w2    s ;s A             Z        �      �      �������c   �������������             ����2    x @x F           Z          �      �      �������c   �������������             ����2    } E} K           �  �        �      �      �������c   �������������             ��2    � J� P           �  v        �      �      �������c   �������������             ,�#�2    � O� U             *        �      �      �������c   �������������             I:�2    � T� Z           J  �        �      �      �������c   �������������             f&Q2    � Y� _           �  �        � 	     �      �������c   �������������         ����    <          d d d d       #   �  �        v        ��        ����c   �������������         ����   " ?          i i i i       %   �  �        v       ��        ����c   �������������         ����   % B          n n n n       '     Z        v       ��        ����c   �������������         ����   ( E          s s s s       )   Z          v       ��       ����c   �������������         ����   + H          x x x x       *   �  �        v       ��       ����c   �������������         ����   . K          } } } }       ,   �  v        v       ��       ����c   �������������         ����   1 N          � � � �       .     *        v       ��       ����c   �������������         ����   4 Q          � � � �       0   J  �        v       ��       ����c   �������������         ����   7 T          � � � �       2   �  �        v       ��       ����c   �������������         ����   : W          � � � �       3   �  F        v	       ��       ����c   �������������         ����     <          d d d d       #   �  �        �        ��        ����c   �������������         ����    " ?          i i i i       %   �  �        �       ��        ����c   �������������         ����    % B          n n n n       '     Z        �       ��        ����c   �������������         ����    ( E          s s s s       )   Z          �       ��       ����c   �������������         ����    + H          x x x x       *   �  �        �       ��       ����c   �������������         ����    . K          } } } }       ,   �  v        �       ��       ����c   �������������         ����    1 N          � � � �       .     *        �       ��       ����c   �������������         ����    4 Q          � � � �       0   J  �        �       ��       ����c   �������������         ����    7 T          � � � �       2   �  �        �       ��       ����c   �������������         ����    : W          � � � �       3   �  F        �	       ��       ����c   �������������         ����� ��                            ����'   N        �      ��i ��        ������  ����������������        ��m ��                         @  S   >C             ��C ��D        ������  ����������������        ��m ��                         `;  Q'  {�             ��D ��E        ������  ����������������        ��m ��                         �Z  /  4             ��E ��F        ������  ����������������        ��m ��                         @�  f7  .�             ��F ��G        ������  ����������������        ��m ��                         �8 }@  ֆ             ��G ��H        ������  ����������������        ��m ��                          q GJ  )Z             ��H ��I        ������  ����������������        ��m ��                    3     ��
 �T  @L             ��I ��J        ������  ����������������        ��m ��                    L     @0 �_  4_             ��J ��K        ������  ����������������        ��m ��                    y     @e �k  �             ��K ��L        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��R ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������        ��t ��                           ����'   N  ?     _      �� ��        ������  ����������������        ��t ��                           ����'   N  ?     `      �� ��        ������  ����������������         ��d ��                          �   �   �        �     ��. ��<        ������  ����������������         ��d ��                          �   �  S        �     ��. ��=        ������  ����������������         ��d ��  (                        �   �  �        �     ��. ��>        ������  ����������������         ��d ��  2                        �   !  �        �     ��. ��?        ������  ����������������         ��e ��                          �   �   �        �     ��/ ��@        ������  ����������������         ��e ��                          �   �  S        �     ��/ ��A        ������  ����������������         ��e ��  (                        �   �  �        �     ��/ ��B        ������  ����������������         ��e ��  2                        �   !  �        �     ��/ ��C        ������  ����������������        ����k ��.1                          ����[
  ">        �      ��; ��        ������  ����������������        ����k ��/1                          �����  �e        �      ��; ��         ������  ����������������        ����k ��01                          ����.  0(       �      ��< ��!        ������  ����������������        ����k ��11                          ����h6  H�       �      ��< ��"        ������  ����������������         ��d ��  P                        �   '  A        �     ��. ��#        ������  ����������������         ��d ��  d                        �   �:  US        �     ��. ��$        ������  ����������������         ��e ��  P                        �   '  A        �     ��/ ��%        ������  ����������������         ��e ��  d                        �   �:  US        �     ��/ ��&        ������  ����������������        ��t ��                           ������  �      a      �� ��        ������  ����������������        ��t ��                           ���� � @B      b      �� ��        ������  ����������������        ��t ��                           ����@B ��      c      �� ��        ������  ����������������        ��} ��    61                    �  '  �� ;     �      �� ��        ������  ����������������        ��} ��                            �  '  ��      �      �� ��        ������  ����������������        ��} ��    >1                       '  �� ;     �      �� ��        ������  ����������������        ��} ��    ?1                    �  '  �� ;     �      �� ��        ������  ����������������        ��} ��    @1                    �I '  �� ;     �      �� ��        ������  ����������������        ��} ��    A1                    �  '  �� ;     �      �� ��        ������  ����������������        ��} ��    B1                    �I '  �� ;     �      �� ��        ������  ����������������        ��} ��    C1                    �O '  �� ;     �      �� ��        ������  ����������������        ��} ��    D1                    �O '  �� ;     �      �� ��        ������  ����������������        ��} ��                               '  ��      �      �� ��        ������  ����������������        ��} ��                            �  '  ��      �      �� ��        ������  ����������������        ��} ��                            �  '  ��      �      �� ��        ������  ����������������        ��} ��                            �I '  ��      �      �� ��        ������  ����������������        ��} ��                            �  '  ��      �      �� ��        ������  ����������������        ��} ��                            �I '  ��      �      �� ��        ������  ����������������        ��} ��                            �O '  ��      �      �� ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������       ����� ��                            ����'   N        �      ��j ��        ������  ����������������          ����E2    ��NB�     ~4  v 8�                  '    ������� � �����  �  �            ���d-2    ��UI�     �4  � ��   ��            '    ������� � �����  �  �            ��-��M2    �\P�     b5  �
 H�   ��            '    ������� � �����  �  �            ��H�m2    �cW�     �5  $ �   ��            '   ������� � �����  �  �            ��c)��2    �j^�     F6  ^ X3   ��            '   ������� � �����  �  �            ��~F��2    �qe�     �6  � �_   ��            '   ������� � �����  �  �            ���c��2    �$xl�     *7  � h�   ��            '   ������� �����  �  �            �����2    �,s�     �7   �   ��            '   ������� 	�����  �  �            ����=	2    4�z�     8  F x�   ��            '   ������� �����  �  �            ����\-	2    <���     �8  �     ��   	         '   �������    �  �  �            ���p�2    � vj�     2=  h# ��   ��             (    ������� � �����  �  �            ����/	2    �(}q�     �=  �% �   ��            (    ������� � �����  �  �            ����P*	2    �0�x�     .>  ( �I   ��            (    ������� � �����  �  �            ����qL	2    8��     �>  p* 0{   ��            (   ������� � �����  �  �            ����n	2    @���     *?  �, h�   ��            (   ������� � �����  �  �            ��)��	2    H���     �?   / ��   ��            (   ������� �����  �  �            ��F$��	2    #P���     &@  x1 �   ��            (   ������� �����  �  �            ��cB��	2    ,X���     �@  �3 @   ��            (   ������� �����  �  �            ���`	�	2    5`���     "A  (6 Hq   ��            (   ������� �����  �  �            ���~7	
2    >h���     �A  �8 ��   ��   	         (   ������� )   �  �  �            ����K2    �NB�     �4  f ��       *       (   )    ������� � �����  �  �            ���d.2    �UI�      5  �	 ��   ��  *      (   )    ������� � �����  �  �            ��=�}I2    �\P�     �5  � �   ��  *      (   )    ������� � �����  �  �            ��^	�d2    �cW�     6   �   ��  *      (   )   ������� � �����  �  �            ��A	�2    �#j^�     v6  N F   ��  *      (   )   ������� � �����  �  �            ���c	��2    �+qe�     �6  � �r   ��  *      (   )   ������� � �����  �  �            ����	��2    �3xl�     Z7  � (�   ��  *      (   )   ������� �����  �  �            ����	��2    ;s�     �7  � ��   ��  *      (   )   ������� 	�����  �  �            ��	�	�2    C�z�     >8  6 8�   ��  *      (   )   ������� �����  �  �            ��$	�	,2    K���     �8  p �$   ��  * 	     (   )   ������� Q   �  �  �            ����	��2    �/vj�     d=  X$ 8�   ��  +       )   *    ������� � �����  �  �            ����	��2    7}q�     �=  �& p,   ��  +      )   *    ������� � �����  �  �            ��	�	�2    ?�x�     `>  ) �]   ��  +      )   *    ������� � �����  �  �            ��A	
)2    G��     �>  `+ ��   ��  +      )   *   ������� � �����  �  �            ��d	6
D*2     O���     \?  �- �   ��  +      )   *   ������� � �����  �  �            ���	Z
_F2    )W���     �?  0 P�   ��  +      )   *   ������� �����  �  �            ���	~
zb2    2_���     X@  h2 �"   ��  +      )   *   ������� �����  �  �            ���	�
�~2    ;g���     �@  �4 �S   ��  +      )   *   ������� �����  �  �            ���	�
��2    Do���     TA  7 ��   ��  +      )   *   ������� �����  �  �            ��
�
��2    Mw���     �A  p9 0�   ��  + 	     )   *   ������� [   �  �  �            ���k�k2    kVkJ�     �4  � �       >       <   +    ������� � �����  �  �            ������2    t]tQ�     �4  � p�   ��  >      <   +    ������� � �����  �  �            ������2    }d}X�     n5  & ��   ��  >      <   +    ������� � �����  �  �            ����2    �k�_�     �5  ` �   ��  >      <   +   ������� � �����  �  �            ��!�!�2    �r�f�     R6  � 8   ��  >      <   +   ������� � �����  �  �            ��>>2    �y�m�     �6  � �d   ��  >      <   +   ������� � �����  �  �            ��[%[%2    ���t�     67   �   ��  >      <   +   ������� �����  �  �            ��xDxD2    ���{�     �7  H ��   ��  >      <   +   ������� 	�����  �  �            ���c�c2    �����     8  � (�   ��  >      <   +   ������� �����  �  �            ������2    �����     �8  � �   ��  > 	     <   +   ������� �   �  �  �            ��b:b:2    �~�r�     >=  �# t�   ��  ?       =   ,    ������� � �����  �  �            ���Z�Z2    ���y�     �=  �% �   ��  ?      =   ,    ������� � �����  �  �            ���z�z2    �����     :>  T( �N   ��  ?      =   ,    ������� � �����  �  �            ������2    �����     �>  �* �   ��  ?      =   ,   ������� � �����  �  �            ������2    �����     6?  - T�   ��  ?      =   ,   ������� � �����  �  �            ������2    �����     �?  \/ ��   ��  ?      =   ,   ������� �����  �  �            ����2    �����     2@  �1 �   ��  ?      =   ,   ������� �����  �  �            ��;	;	2    �����     �@  4 �D   ��  ?      =   ,   ������� �����  �  �            ��Z:	Z:	2    �����     .A  d6 4v   ��  ?      =   ,   ������� �����  �  �            ��yZ	yZ	2    �����     �A  �8 l�   ��  ? 	     =   ,   ������� �   �  �  �            ��E��2    ��NB�     �4  * H�       T       Q   -    ������� � �����  �  �            ��d-�2    �UI�     5  d	 л   ��  T      Q   -    ������� � �����  �  �            ���M-�2    �\P�     �5  � X�   ��  T      Q   -    ������� � �����  �  �            ���mH2    �cW�     �5  � �   ��  T      Q   -   ������� � �����  �  �            ����c)2    �j^�     j6   hA   ��  T      Q   -   ������� � �����  �  �            ����~F2    �&qe�     �6  L �m   ��  T      Q   -   ������� � �����  �  �            �����c2    �.xl�     N7  � x�   ��  T      Q   -   ������� �����  �  �            �����2    6s�     �7  �  �   ��  T      Q   -   ������� 	�����  �  �            ��=	��2    >�z�     28  � ��   ��  T      Q   -   ������� �����  �  �            ��\-	��2    F���     �8  4     ��  T 	     Q   -   ������� �   �  �  �            ����p2    �*vj�     W=  $ L�   ��  U       R   .    ������� � �����  �  �            ��/	��2     2}q�     �=  t& �'   ��  U      R   .    ������� � �����  �  �            ��P*	��2    	:�x�     S>  �( �X   ��  U      R   .    ������� � �����  �  �            ��qL	��2    B��     �>  $+ �   ��  U      R   .   ������� � �����  �  �            ���n	�2    J���     O?  |- ,�   ��  U      R   .   ������� � �����  �  �            ����	)2    $R���     �?  �/ d�   ��  U      R   .   ������� �����  �  �            ����	F$2    -Z���     K@  ,2 �   ��  U      R   .   ������� �����  �  �            ����	cB2    6b���     �@  �4 �N   ��  U      R   .   ������� �����  �  �            ��	�	�`2    ?j���     GA  �6 �   ��  U      R   .   ������� �����  �  �            ��7	
�~2    Hr���     �A  49 D�   ��  U 	     R   .   ������� �   �  �  �            ��K��2    s��H�     r4  : �|       j       f   /    ������� � �����  �  �            ��d.�2    z��O�     �4  t �   ��  j      f   /    ������� � �����  �  �            ��}I=�2    ���V�     V5  �
 ��   ��  j      f   /    ������� � �����  �  �            ���d^	2    ���]�     �5  �     ��  j      f   /   ������� � �����  �  �            ���A	2    ���d�     :6  " �.   ��  j      f   /   ������� � �����  �  �            �����c	2    ���k�     �6  \ 0[   ��  j      f   /   ������� � �����  �  �            ������	2    � �r�     7  � ��   ��  j      f   /   ������� �����  �  �            ������	2    ��y�     �7  � @�   ��  j      f   /   ������� 	�����  �  �            ���	�	2    ���     8  
 ��   ��  j      f   /   ������� �����  �  �            ��,$	�	2    ���     t8  D P   ��  j 	     f   /   ������� �   �  �  �            ������	2    ���p�     %=  ,# ��   ��  k       g   0    ������� � �����  �  �            ������	2    ��w�     �=  �% �   ��  k      g   0    ������� � �����  �  �            ���	�	2    �~�     !>  �' E   ��  k      g   0    ������� � �����  �  �            ��)A	
2    ���     �>  4* Dv   ��  k      g   0   ������� � �����  �  �            ��D*d	6
2    ���     ?  �, |�   ��  k      g   0   ������� � �����  �  �            ��_F�	Z
2    �&��     �?  �. ��   ��  k      g   0   ������� �����  �  �            ��zb�	~
2    �.(��     @  <1 �	   ��  k      g   0   ������� �����  �  �            ���~�	�
2    �61��     �@  �3 $;   ��  k      g   0   ������� �����  �  �            �����	�
2    �>:��     A  �5 \l   ��  k      g   0   ������� �����  �  �            ����
�
2    �FC��     �A  D8 ��   ��  k 	     g   0   ������� �   �  �  �             HH
2    iVkJ�     �4  � ��       �       ~   1    ������� � �����  �  �             d$d$
2    r]tQ�     5  (	  �   ��  �      ~   1    ������� � �����  �  �             �B�B
2    {d}X�     z5  b ��   ��  �      ~   1    ������� � �����  �  �             �`�`
2    �k�_�     �5  � 0   ��  �      ~   1   ������� � �����  �  �             �~�~
2    �r�f�     ^6  � �<   ��  �      ~   1   ������� � �����  �  �             ����
2    �y�m�     �6   @i   ��  �      ~   1   ������� � �����  �  �             ����
2    ���t�     B7  J ȕ   ��  �      ~   1   ������� �����  �  �             ��
2    ���{�     �7  � P�   ��  �      ~   1   ������� 	�����  �  �             (�(�
2    �����     &8  � ��   ��  �      ~   1   ������� �����  �  �             DD
2    �����     �8  � `   ��  � 	     ~   1   �������   �  �  �             ����
2    �~�r�     K=  �# `�   ��  �          2    ������� � �����  �  �             ��
2    ���y�     �=  8& �"   ��  �         2    ������� � �����  �  �             /	/	
2    �����     G>  �( �S   ��  �         2    ������� � �����  �  �             M(M(
2    �����     �>  �* �   ��  �         2   ������� � �����  �  �             kGkG
2    �����     C?  @- @�   ��  �         2   ������� � �����  �  �             �f�f
2    �����     �?  �/ x�   ��  �         2   ������� �����  �  �             ����
2    �����     ?@  �1 �   ��  �         2   ������� �����  �  �             ����
2    �����     �@  H4 �I   ��  �         2   ������� �����  �  �             ����
2    �����     ;A  �6  {   ��  �         2   ������� �����  �  �             ��
2    �����     �A  �8 X�   ��  � 	        2   ������� #  �  �  �             �lK2    �NB�     �4  f ��       �       �   3    ������� � �����  �  �             ��d.2    �UI�      5  �	 ��   ��  �      �   3    ������� � �����  �  �             ��}I2    !�\P�     �5  � �   ��  �      �   3    ������� � �����  �  �             ���d2    )�cW�     6   �   ��  �      �   3   ������� � �����  �  �             ��2    1�j^�     v6  N F   ��  �      �   3   ������� � �����  �  �             0	��2    9�qe�     �6  � �r   ��  �      �   3   ������� � �����  �  �             P2	��2    A�xl�     Z7  � (�   ��  �      �   3   ������� �����  �  �             pS	��2    I�s�     �7  � ��   ��  �      �   3   ������� 	�����  �  �             �t	�2    Q��z�     >8  6 8�   ��  �      �   3   ������� �����  �  �             ��	,2    Y����     �8  p �$   ��  � 	     �   3   �������    �  �  �             cO	��2    <�vj�     d=  X$ 8�   ��  �       �   4    ������� � �����  �  �             �r	��2    D�}q�     �=  �& p,   ��  �      �   4    ������� � �����  �  �             ��	�2    L��x�     `>  ) �]   ��  �      �   4    ������� � �����  �  �             ��	)2    T���     �>  `+ ��   ��  �      �   4   ������� � �����  �  �             ��	D*2    \����     \?  �- �   ��  �      �   4   ������� � �����  �  �             	�	_F2    d����     �?  0 P�   ��  �      �   4   ������� �����  �  �             /	!
zb2    l����     X@  h2 �"   ��  �      �   4   ������� �����  �  �             Q	D
�~2    t���     �@  �4 �S   ��  �      �   4   ������� �����  �  �             s	g
��2    |���     TA  7 ��   ��  �      �   4   ������� �����  �  �             �	�
��2    ����     �A  p9 0�   ��  � 	     �   4   ������� )   �  �  �         ����   F G          5� � �     C    ^N   ��  #        ��5        ���� �����  �  �         ����   H I          <� � �     �  f�  �f   ��  #       ��5        ���� �����  �  �         ����   J K          C� � �     �  
�  �   ��  #       ��5        ���� �����  �  �         ����   M N          J� � �        ��  2�   ��  #       ��5       ���� �����  �  �         ����   O P          %Q� � �     ?  R�  ΰ   ��  #       ��5       ���� �����  �  �         ����   Q R          -X� � �     ~  ��  j�   ��  #       ��5       ���� �����  �  �         ����   S T          5_� � �     �  ��  �   ��  #       ��5       ���� �����  �  �         ����   U V          =f� � �     �  >�  ��   ��  #       ��5       ���� �����  �  �         ����   X Y          Em� � �     ;  �  >	   ��  #       ��5       ���� &�����  �  �         ����   Z [          Mt� � �     z  ��  �+	   ��  #	       ��5       ���� /K  �  �  �         ����   K L          3[� � �       �  `1
   ��  $        ��6        ���� �����  �  �         ����   M N          ;b� � �     `  ؤ  �M
   ��  $       ��6        ���� �����  �  �         ����   O P          Ci� � �     �  ��  �i
   ��  $       ��6        ���� �����  �  �         ����   R S          Kp� � �     �  \�  ��
   ��  $       ��6       ���� �����  �  �         ����   T U          Sw� � �     8  �  �
   ��  $       ��6       ���� �����  �  �         ����   V W          [~� � �     �  �   �
   ��  $       ��6       ���� �����  �  �         ����   X Y          c�� � �     �  ��   �
   ��  $       ��6       ���� $�����  �  �         ����   Z [          k�� � �       d�  @�
   ��  $       ��6       ���� +�����  �  �         ����   ] ^          s�� �     X  &�  `   ��  $       ��6       ���� 3�����  �  �         ����   _ `          {�� �     �  �  �.   ��  $	       ��6       ���� <U  �  �  �         ����   7 8          � 3�� �     C    ^N   ��  7        ��7        ���� �����  �  �         ����   9 :          � 9� �     �  f�  �f   ��  7       ��7        ���� �����  �  �         ����   ; <          � ?� �     �  
�  �   ��  7       ��7        ���� �����  �  �         ����   = >          � E� �        ��  2�   ��  7       ��7       ���� �����  �  �         ����   ? @          � K� �     ?  R�  ΰ   ��  7       ��7       ���� �����  �  �         ����   A B          Q&� �     ~  ��  j�   ��  7       ��7       ���� �����  �  �         ����   D E          W.� �     �  ��  �   ��  7       ��7       ���� �����  �  �         ����   F G          ]6� �     �  >�  ��   ��  7       ��7       ���� �����  �  �         ����   H I          c>� �     ;  �  >	   ��  7       ��7       ���� &�����  �  �         ����   J K          iF� �     z  ��  �+	   ��  7	       ��7       ���� /K  �  �  �         ����   ; <          P,� �       �  `1
   ��  8        ��8        ���� �����  �  �         ����   = >          
W4� �     `  ؤ  �M
   ��  8       ��8        ���� �����  �  �         ����   ? @          ^<� �     �  ��  �i
   ��  8       ��8        ���� �����  �  �         ����   A B          eD� �     �  \�  ��
   ��  8       ��8       ���� �����  �  �         ����   C D          lL� �     8  �  �
   ��  8       ��8       ���� �����  �  �         ����   E F          "sT� �     �  �   �
   ��  8       ��8       ���� �����  �  �         ����   H I          (z\� �     �  ��   �
   ��  8       ��8       ���� $�����  �  �         ����   J K          .�d� �       d�  @�
   ��  8       ��8       ���� +�����  �  �         ����   L M          4�l� �     X  &�  `   ��  8       ��8       ���� 3�����  �  �         ����   N O          :�t�     �  �  �.   ��  8	       ��8       ���� <U  �  �  �         ����   6 7          �� �� �     C    ^N   ��  K        ��9        ���� �����  �  �         ����   8 9          �� �� �     �  f�  �f   ��  K       ��9        ���� �����  �  �         ����   : ;          �� �� �     �  
�  �   ��  K       ��9        ���� �����  �  �         ����   < =          �� �� �        ��  2�   ��  K       ��9       ���� �����  �  �         ����   > ?          �� �� �     ?  R�  ΰ   ��  K       ��9       ���� �����  �  �         ����   @ A          �� �� �     ~  ��  j�   ��  K       ��9       ���� �����  �  �         ����   C D          �� �� �     �  ��  �   ��  K       ��9       ���� �����  �  �         ����   E F          �� �� �     �  >�  ��   ��  K       ��9       ���� �����  �  �         ����   G H          �� �� �     ;  �  >	   ��  K       ��9       ���� &�����  �  �         ����   I J          �� �� �     z  ��  �+	   ��  K	       ��9       ���� /K  �  �  �         ����   : ;          �� �� �       �  `1
   ��  L        ��:        ���� �����  �  �         ����   < =          �� �� �     `  ؤ  �M
   ��  L       ��:        ���� �����  �  �         ����   > ?          �� �� �     �  ��  �i
   ��  L       ��:        ���� �����  �  �         ����   @ A          �� �� �     �  \�  ��
   ��  L       ��:       ���� �����  �  �         ����   B C          �� �� �     8  �  �
   ��  L       ��:       ���� �����  �  �         ����   D E          �� �� �     �  �   �
   ��  L       ��:       ���� �����  �  �         ����   G H          � � �     �  ��   �
   ��  L       ��:       ���� $�����  �  �         ����   I J          	� 	� �       d�  @�
   ��  L       ��:       ���� +�����  �  �         ����   K L          � � �     X  &�  `   ��  L       ��:       ���� 3�����  �  �         ����   M N          � � �     �  �  �.   ��  L	       ��:       ���� <U  �  �  �         ����   ) *          � ( � �     C    ^N   ��  _        ��;        ���� �����  �  �         ����   + ,          � .� �     �  f�  �f   ��  _       ��;        ���� �����  �  �         ����   - .          � 4� �     �  
�  �   ��  _       ��;        ���� �����  �  �         ����   / 0          � :� �        ��  2�   ��  _       ��;       ���� �����  �  �         ����   1 2          � @ � �     ?  R�  ΰ   ��  _       ��;       ���� �����  �  �         ����   3 4          � F(� �     ~  ��  j�   ��  _       ��;       ���� �����  �  �         ����   5 6          � L0� �     �  ��  �   ��  _       ��;       ���� �����  �  �         ����   7 8          � R8� �     �  >�  ��   ��  _       ��;       ���� �����  �  �         ����   9 :          � X@� �     ;  �  >	   ��  _       ��;       ���� &�����  �  �         ����   ; <          ^H� �     z  ��  �+	   ��  _	       ��;       ���� /K  �  �  �         ����   , -          � E.� �       �  `1
   ��  `        ��<        ���� �����  �  �         ����   . /          � L6� �     `  ؤ  �M
   ��  `       ��<        ���� �����  �  �         ����   0 1          � S>� �     �  ��  �i
   ��  `       ��<        ���� �����  �  �         ����   2 3          ZF� �     �  \�  ��
   ��  `       ��<       ���� �����  �  �         ����   4 5          aN� �     8  �  �
   ��  `       ��<       ���� �����  �  �         ����   6 7          hV� �     �  �   �
   ��  `       ��<       ���� �����  �  �         ����   8 9          o^� �     �  ��   �
   ��  `       ��<       ���� $�����  �  �         ����   : ;          vf� �       d�  @�
   ��  `       ��<       ���� +�����  �  �         ����   < =          }n� �     X  &�  `   ��  `       ��<       ���� 3�����  �  �         ����   > ?          %�v�     �  �  �.   ��  `	       ��<       ���� <U  �  �  �         ����   7 8          ��� � �     C    ^N   ��  s        ��=        ���� �����  �  �         ����   9 :          ��� � �     �  f�  �f   ��  s       ��=        ���� �����  �  �         ����   ; <          ��� � �     �  
�  �   ��  s       ��=        ���� �����  �  �         ����   = >          ��� � �        ��  2�   ��  s       ��=       ���� �����  �  �         ����   ? @          ��� � �     ?  R�  ΰ   ��  s       ��=       ���� �����  �  �         ����   A B          ��� � �     ~  ��  j�   ��  s       ��=       ���� �����  �  �         ����   D E          ��� � �     �  ��  �   ��  s       ��=       ���� �����  �  �         ����   F G          ��� � �     �  >�  ��   ��  s       ��=       ���� �����  �  �         ����   H I          ��� � �     ;  �  >	   ��  s       ��=       ���� &�����  �  �         ����   J K          ��� � �     z  ��  �+	   ��  s	       ��=       ���� /K  �  �  �         ����   ; <          ��� � �       �  `1
   ��  t        ��>        ���� �����  �  �         ����   = >          ��� � �     `  ؤ  �M
   ��  t       ��>        ���� �����  �  �         ����   ? @          ��� � �     �  ��  �i
   ��  t       ��>        ���� �����  �  �         ����   A B          ��� � �     �  \�  ��
   ��  t       ��>       ���� �����  �  �         ����   C D          ��� � �     8  �  �
   ��  t       ��>       ���� �����  �  �         ����   E F          ��� � �     �  �   �
   ��  t       ��>       ���� �����  �  �         ����   H I          ��� � �     �  ��   �
   ��  t       ��>       ���� $�����  �  �         ����   J K          ��� � �       d�  @�
   ��  t       ��>       ���� +�����  �  �         ����   L M          ��� �     X  &�  `   ��  t       ��>       ���� 3�����  �  �         ����   N O          ��� �     �  �  �.   ��  t	       ��>       ���� <U  �  �  �         ����    6 7          � !�� �     C    ^N   ��  �        ��?        ���� �����  �  �         ����    8 9          � ' � �     �  f�  �f   ��  �       ��?        ���� �����  �  �         ����    : ;          � -� �     �  
�  �   ��  �       ��?        ���� �����  �  �         ����    < =          � 3� �        ��  2�   ��  �       ��?       ���� �����  �  �         ����    > ?          � 9� �     ?  R�  ΰ   ��  �       ��?       ���� �����  �  �         ����    @ A          � ? � �     ~  ��  j�   ��  �       ��?       ���� �����  �  �         ����    C D          � E(� �     �  ��  �   ��  �       ��?       ���� �����  �  �         ����    E F          � K0� �     �  >�  ��   ��  �       ��?       ���� �����  �  �         ����    G H           Q8� �     ;  �  >	   ��  �       ��?       ���� &�����  �  �         ����    I J          W@� �     z  ��  �+	   ��  �	       ��?       ���� /K  �  �  �         ����    : ;          � >&� �       �  `1
   ��  �        ��@        ���� �����  �  �         ����    < =          � E.� �     `  ؤ  �M
   ��  �       ��@        ���� �����  �  �         ����    > ?          � L6� �     �  ��  �i
   ��  �       ��@        ���� �����  �  �         ����    @ A          S>� �     �  \�  ��
   ��  �       ��@       ���� �����  �  �         ����    B C          ZF� �     8  �  �
   ��  �       ��@       ���� �����  �  �         ����    D E          aN� �     �  �   �
   ��  �       ��@       ���� �����  �  �         ����    G H          hV� �     �  ��   �
   ��  �       ��@       ���� $�����  �  �         ����    I J          o^� �       d�  @�
   ��  �       ��@       ���� +�����  �  �         ����    K L           vf� �     X  &�  `   ��  �       ��@       ���� 3�����  �  �         ����    M N          &}n� �     �  �  �.   ��  �	       ��@       ���� <U  �  �  �         ����  D E          �5� � �     �  ΋  1   ��  �        ��A        ���� �����  �  �         ����  F G          �<� � �     7  r�  �I   ��  �       ��A        ���� �����  �  �         ����  H I           C� � �     v  �  Jb   ��  �       ��A        ���� �����  �  �         ����  K L          J� � �     �  ��  �z   ��  �       ��A       ���� �����  �  �         ����  M N          Q� � �     �  ^�  ��   ��  �       ��A       ���� �����  �  �         ����  O P          X� � �     3  �  �   ��  �       ��A       ���� �����  �  �         ����  Q R           _� � �     r  ��  ��   ��  �       ��A       ���� �����  �  �         ����  S T          (f� � �     �  J�  V�   ��  �       ��A       ���� �����  �  �         ����  V W          0m� � �     �  �  ��   ��  �       ��A       ���� &�����  �  �         ����  X Y          8t� � �     /  ��  �	   ��  �	       ��A       ���� /K  �  �  �         ����  I J          [� � �     �  "�   
   ��  �        ��B        ���� �����  �  �         ����  K L          &b� � �       �  @.
   ��  �       ��B        ���� �����  �  �         ����  M N          .i� � �     X  ��  `J
   ��  �       ��B        ���� �����  �  �         ����  P Q          6p� � �     �  h�  �f
   ��  �       ��B       ���� �����  �  �         ����  R S          >w� � �     �  *�  ��
   ��  �       ��B       ���� �����  �  �         ����  T U          F~� � �     0  �  ��
   ��  �       ��B       ���� �����  �  �         ����  V W          N�� � �     x  ��  �
   ��  �       ��B       ���� $�����  �  �         ����  X Y          V�� � �     �  p�   �
   ��  �       ��B       ���� +�����  �  �         ����  [ \          ^�� �       2�   �
   ��  �       ��B       ���� 3�����  �  �         ����  ] ^          f�� �     P  ��  @   ��  �	       ��B       ���� <U  �  �  �         ����  6 7          � �� �     �  ΋  1   ��  �        ��C        ���� �����  �  �         ����  8 9          � $�� �     7  r�  �I   ��  �       ��C        ���� �����  �  �         ����  : ;          � *�� �     v  �  Jb   ��  �       ��C        ���� �����  �  �         ����  < =          � 0� �     �  ��  �z   ��  �       ��C       ���� �����  �  �         ����  > ?          � 6	� �     �  ^�  ��   ��  �       ��C       ���� �����  �  �         ����  @ A          � <� �     3  �  �   ��  �       ��C       ���� �����  �  �         ����  C D          � B� �     r  ��  ��   ��  �       ��C       ���� �����  �  �         ����  E F          � H!� �     �  J�  V�   ��  �       ��C       ���� �����  �  �         ����  G H          � N)� �     �  �  ��   ��  �       ��C       ���� &�����  �  �         ����  I J          T1� �     /  ��  �	   ��  �	       ��C       ���� /K  �  �  �         ����  : ;          � ;� �     �  "�   
   ��  �        ��D        ���� �����  �  �         ����  < =          � B� �       �  @.
   ��  �       ��D        ���� �����  �  �         ����  > ?          � I'� �     X  ��  `J
   ��  �       ��D        ���� �����  �  �         ����  @ A          P/� �     �  h�  �f
   ��  �       ��D       ���� �����  �  �         ����  B C          W7� �     �  *�  ��
   ��  �       ��D       ���� �����  �  �         ����  D E          ^?� �     0  �  ��
   ��  �       ��D       ���� �����  �  �         ����  G H          eG� �     x  ��  �
   ��  �       ��D       ���� $�����  �  �         ����  I J          lO� �     �  p�   �
   ��  �       ��D       ���� +�����  �  �         ����  K L          sW� �       2�   �
   ��  �       ��D       ���� 3�����  �  �         ����  M N          %z_�     P  ��  @   ��  �	       ��D       ���� <U  �  �  �         ����  5 6          �� �� �     �  ΋  1   ��  �        ��E        ���� �����  �  �         ����  7 8          �� �� �     7  r�  �I   ��  �       ��E        ���� �����  �  �         ����  9 :          �� �� �     v  �  Jb   ��  �       ��E        ���� �����  �  �         ����  ; <          �� �� �     �  ��  �z   ��  �       ��E       ���� �����  �  �         ����  = >          �� �� �     �  ^�  ��   ��  �       ��E       ���� �����  �  �         ����  ? @          �� �� �     3  �  �   ��  �       ��E       ���� �����  �  �         ����  B C          �� �� �     r  ��  ��   ��  �       ��E       ���� �����  �  �         ����  D E          �� �� �     �  J�  V�   ��  �       ��E       ���� �����  �  �         ����  F G          �� �� �     �  �  ��   ��  �       ��E       ���� &�����  �  �         ����  H I          �� �� �     /  ��  �	   ��  �	       ��E       ���� /K  �  �  �         ����  9 :          �� �� �     �  "�   
   ��  �        ��F        ���� �����  �  �         ����  ; <          �� �� �       �  @.
   ��  �       ��F        ���� �����  �  �         ����  = >          �� �� �     X  ��  `J
   ��  �       ��F        ���� �����  �  �         ����  ? @          �� �� �     �  h�  �f
   ��  �       ��F       ���� �����  �  �         ����  A B          �� �� �     �  *�  ��
   ��  �       ��F       ���� �����  �  �         ����  C D          �� �� �     0  �  ��
   ��  �       ��F       ���� �����  �  �         ����  F G          �� �� �     x  ��  �
   ��  �       ��F       ���� $�����  �  �         ����  H I          �� �� �     �  p�   �
   ��  �       ��F       ���� +�����  �  �         ����  J K          �� �� �       2�   �
   ��  �       ��F       ���� 3�����  �  �         ����  L M          � � �     P  ��  @   ��  �	       ��F       ���� <U  �  �  �         ����  ( )          � �� �     �  ΋  1   ��  �        ��G        ���� �����  �  �         ����  * +          � %�� �     7  r�  �I   ��  �       ��G        ���� �����  �  �         ����  , -          � +� �     v  �  Jb   ��  �       ��G        ���� �����  �  �         ����  . /          � 1� �     �  ��  �z   ��  �       ��G       ���� �����  �  �         ����  0 1          � 7� �     �  ^�  ��   ��  �       ��G       ���� �����  �  �         ����  2 3          � =� �     3  �  �   ��  �       ��G       ���� �����  �  �         ����  4 5          � C'� �     r  ��  ��   ��  �       ��G       ���� �����  �  �         ����  6 7          � I/� �     �  J�  V�   ��  �       ��G       ���� �����  �  �         ����  8 9          � O7� �     �  �  ��   ��  �       ��G       ���� &�����  �  �         ����  : ;          � U?� �     /  ��  �	   ��  �	       ��G       ���� /K  �  �  �         ����  + ,          � <%� �     �  "�   
   ��  �        ��H        ���� �����  �  �         ����  - .          � C-� �       �  @.
   ��  �       ��H        ���� �����  �  �         ����  / 0          � J5� �     X  ��  `J
   ��  �       ��H        ���� �����  �  �         ����  1 2          � Q=� �     �  h�  �f
   ��  �       ��H       ���� �����  �  �         ����  3 4          � XE� �     �  *�  ��
   ��  �       ��H       ���� �����  �  �         ����  5 6          _M� �     0  �  ��
   ��  �       ��H       ���� �����  �  �         ����  7 8          
fU� �     x  ��  �
   ��  �       ��H       ���� $�����  �  �         ����  9 :          m]� �     �  p�   �
   ��  �       ��H       ���� +�����  �  �         ����  ; <          te� �       2�   �
   ��  �       ��H       ���� 3�����  �  �         ����  = >          {m� �     P  ��  @   ��  �	       ��H       ���� <U  �  �  �         ����  7 8          ��� � �     �  ΋  1   ��  �        ��I        ���� �����  �  �         ����  9 :          ��� � �     7  r�  �I   ��  �       ��I        ���� �����  �  �         ����  ; <          ��� � �     v  �  Jb   ��  �       ��I        ���� �����  �  �         ����  = >          ��� � �     �  ��  �z   ��  �       ��I       ���� �����  �  �         ����  ? @          ��� � �     �  ^�  ��   ��  �       ��I       ���� �����  �  �         ����  A B          ��� � �     3  �  �   ��  �       ��I       ���� �����  �  �         ����  D E          ��� � �     r  ��  ��   ��  �       ��I       ���� �����  �  �         ����  F G          ��� � �     �  J�  V�   ��  �       ��I       ���� �����  �  �         ����  H I          ��� � �     �  �  ��   ��  �       ��I       ���� &�����  �  �         ����  J K          ��� � �     /  ��  �	   ��  �	       ��I       ���� /K  �  �  �         ����  ; <          ��� � �     �  "�   
   ��  �        ��J        ���� �����  �  �         ����  = >          ��� � �       �  @.
   ��  �       ��J        ���� �����  �  �         ����  ? @          ��� � �     X  ��  `J
   ��  �       ��J        ���� �����  �  �         ����  A B          ��� � �     �  h�  �f
   ��  �       ��J       ���� �����  �  �         ����  C D          ��� � �     �  *�  ��
   ��  �       ��J       ���� �����  �  �         ����  E F          ��� � �     0  �  ��
   ��  �       ��J       ���� �����  �  �         ����  H I          ��� � �     x  ��  �
   ��  �       ��J       ���� $�����  �  �         ����  J K          ��� � �     �  p�   �
   ��  �       ��J       ���� +�����  �  �         ����  L M          ��� �       2�   �
   ��  �       ��J       ���� 3�����  �  �         ����  N O          ��� �     P  ��  @   ��  �	       ��J       ���� <U  �  �  �         ����   5 6          � !�� �     �  ΋  1   ��  �        ��K        ���� �����  �  �         ����   7 8          � '�� �     7  r�  �I   ��  �       ��K        ���� �����  �  �         ����   9 :          � -�� �     v  �  Jb   ��  �       ��K        ���� �����  �  �         ����   ; <          � 3� �     �  ��  �z   ��  �       ��K       ���� �����  �  �         ����   = >          � 9� �     �  ^�  ��   ��  �       ��K       ���� �����  �  �         ����   ? @          � ?� �     3  �  �   ��  �       ��K       ���� �����  �  �         ����   B C          � E� �     r  ��  ��   ��  �       ��K       ���� �����  �  �         ����   D E          � K$� �     �  J�  V�   ��  �       ��K       ���� �����  �  �         ����   F G           Q,� �     �  �  ��   ��  �       ��K       ���� &�����  �  �         ����   H I          W4� �     /  ��  �	   ��  �	       ��K       ���� /K  �  �  �         ����   9 :          � >� �     �  "�   
   ��  �        ��L        ���� �����  �  �         ����   ; <          � E"� �       �  @.
   ��  �       ��L        ���� �����  �  �         ����   = >          � L*� �     X  ��  `J
   ��  �       ��L        ���� �����  �  �         ����   ? @          S2� �     �  h�  �f
   ��  �       ��L       ���� �����  �  �         ����   A B          Z:� �     �  *�  ��
   ��  �       ��L       ���� �����  �  �         ����   C D          aB� �     0  �  ��
   ��  �       ��L       ���� �����  �  �         ����   F G          hJ� �     x  ��  �
   ��  �       ��L       ���� $�����  �  �         ����   H I          oR� �     �  p�   �
   ��  �       ��L       ���� +�����  �  �         ����   J K           vZ� �       2�   �
   ��  �       ��L       ���� 3�����  �  �         ����   L M          &}b� �     P  ��  @   ��  �	       ��L       ���� <U  �  �  �         ����  E F          �5� � �     �  j�  6+   ��  �        ��M        ���� �����  �  �         ����  G H          <� � �     (  �  �C   ��  �       ��M        ���� �����  �  �         ����  I J          C� � �     g  ��  n\   ��  �       ��M        ���� �����  �  �         ����  L M          J� � �     �  V�  
u   ��  �       ��M       ���� �����  �  �         ����  N O          Q� � �     �  ��  ��   ��  �       ��M       ���� �����  �  �         ����  P Q          %X� � �     $  ��  B�   ��  �       ��M       ���� �����  �  �         ����  R S          -_� � �     c  B�  ޾   ��  �       ��M       ���� �����  �  �         ����  T U          5f� � �     �  �  z�   ��  �       ��M       ���� �����  �  �         ����  W X          =m� � �     �  ��  �   ��  �       ��M       ���� &�����  �  �         ����  Y Z          Et� � �        .�  �	   ��  �	       ��M       ���� /K  �  �  �         ����  J K          +[� � �     �  ��  �
   ��  �        ��N        ���� �����  �  �         ����  L M          3b� � �        ��   (
   ��  �       ��N        ���� �����  �  �         ����  N O          ;i� � �     H  B�   D
   ��  �       ��N        ���� �����  �  �         ����  Q R          Cp� � �     �  �  @`
   ��  �       ��N       ���� �����  �  �         ����  S T          Kw� � �     �  Ƨ  `|
   ��  �       ��N       ���� �����  �  �         ����  U V          S~� � �        ��  ��
   ��  �       ��N       ���� �����  �  �         ����  W X          [�� � �     h  J�  ��
   ��  �       ��N       ���� $�����  �  �         ����  Y Z          c�� � �     �  �  ��
   ��  �       ��N       ���� +�����  �  �         ����  \ ]          k�� �     �  ή  ��
   ��  �       ��N       ���� 3�����  �  �         ����  ^ _          s�� �     @  ��   	   ��  �	       ��N       ���� <U  �  �  �         ����  6 7          � +�� �     �  j�  6+   ��          ��O        ���� �����  �  �         ����  8 9          � 1�� �     (  �  �C   ��         ��O        ���� �����  �  �         ����  : ;          � 7� �     g  ��  n\   ��         ��O        ���� �����  �  �         ����  < =          � =� �     �  V�  
u   ��         ��O       ���� �����  �  �         ����  > ?          � C� �     �  ��  ��   ��         ��O       ���� �����  �  �         ����  @ A          � I� �     $  ��  B�   ��         ��O       ���� �����  �  �         ����  C D           O&� �     c  B�  ޾   ��         ��O       ���� �����  �  �         ����  E F          U.� �     �  �  z�   ��         ��O       ���� �����  �  �         ����  G H          [6� �     �  ��  �   ��         ��O       ���� &�����  �  �         ����  I J          a>� �        .�  �	   ��  	       ��O       ���� /K  �  �  �         ����  : ;          � H$� �     �  ��  �
   ��          ��P        ���� �����  �  �         ����  < =          O,� �        ��   (
   ��         ��P        ���� �����  �  �         ����  > ?          V4� �     H  B�   D
   ��         ��P        ���� �����  �  �         ����  @ A          ]<� �     �  �  @`
   ��         ��P       ���� �����  �  �         ����  B C          dD� �     �  Ƨ  `|
   ��         ��P       ���� �����  �  �         ����  D E          kL� �        ��  ��
   ��         ��P       ���� �����  �  �         ����  G H           rT� �     h  J�  ��
   ��         ��P       ���� $�����  �  �         ����  I J          &y\� �     �  �  ��
   ��         ��P       ���� +�����  �  �         ����  K L          ,�d� �     �  ή  ��
   ��         ��P       ���� 3�����  �  �         ����  M N          2�l�     @  ��   	   ��  	       ��P       ���� <U  �  �  �         ����  5 6          �� �� �     �  j�  6+   ��          ��Q        ���� �����  �  �         ����  7 8          �� �� �     (  �  �C   ��         ��Q        ���� �����  �  �         ����  9 :          �� �� �     g  ��  n\   ��         ��Q        ���� �����  �  �         ����  ; <          �� �� �     �  V�  
u   ��         ��Q       ���� �����  �  �         ����  = >          �� �� �     �  ��  ��   ��         ��Q       ���� �����  �  �         ����  ? @          �� �� �     $  ��  B�   ��         ��Q       ���� �����  �  �         ����  B C          �� �� �     c  B�  ޾   ��         ��Q       ���� �����  �  �         ����  D E          �� �� �     �  �  z�   ��         ��Q       ���� �����  �  �         ����  F G          �� �� �     �  ��  �   ��         ��Q       ���� &�����  �  �         ����  H I          �� �� �        .�  �	   ��  	       ��Q       ���� /K  �  �  �         ����  9 :          �� �� �     �  ��  �
   ��           ��R        ���� �����  �  �         ����  ; <          �� �� �        ��   (
   ��          ��R        ���� �����  �  �         ����  = >          �� �� �     H  B�   D
   ��          ��R        ���� �����  �  �         ����  ? @          �� �� �     �  �  @`
   ��          ��R       ���� �����  �  �         ����  A B          �� �� �     �  Ƨ  `|
   ��          ��R       ���� �����  �  �         ����  C D          �� �� �        ��  ��
   ��          ��R       ���� �����  �  �         ����  F G          �� �� �     h  J�  ��
   ��          ��R       ���� $�����  �  �         ����  H I          � � �     �  �  ��
   ��          ��R       ���� +�����  �  �         ����  J K          	� 	� �     �  ή  ��
   ��          ��R       ���� 3�����  �  �         ����  L M          � � �     @  ��   	   ��   	       ��R       ���� <U  �  �  �         ����  ( )          � *�� �     �  j�  6+   ��  0        ��S        ���� �����  �  �         ����  * +          � 0� �     (  �  �C   ��  0       ��S        ���� �����  �  �         ����  , -          � 6
� �     g  ��  n\   ��  0       ��S        ���� �����  �  �         ����  . /          � <� �     �  V�  
u   ��  0       ��S       ���� �����  �  �         ����  0 1          � B� �     �  ��  ��   ��  0       ��S       ���� �����  �  �         ����  2 3          � H"� �     $  ��  B�   ��  0       ��S       ���� �����  �  �         ����  4 5          � N*� �     c  B�  ޾   ��  0       ��S       ���� �����  �  �         ����  6 7          T2� �     �  �  z�   ��  0       ��S       ���� �����  �  �         ����  8 9          Z:� �     �  ��  �   ��  0       ��S       ���� &�����  �  �         ����  : ;          `B� �        .�  �	   ��  0	       ��S       ���� /K  �  �  �         ����  + ,          � G(� �     �  ��  �
   ��  1        ��T        ���� �����  �  �         ����  - .          � N0� �        ��   (
   ��  1       ��T        ���� �����  �  �         ����  / 0          U8� �     H  B�   D
   ��  1       ��T        ���� �����  �  �         ����  1 2          
\@� �     �  �  @`
   ��  1       ��T       ���� �����  �  �         ����  3 4          cH� �     �  Ƨ  `|
   ��  1       ��T       ���� �����  �  �         ����  5 6          jP� �        ��  ��
   ��  1       ��T       ���� �����  �  �         ����  7 8          qX� �     h  J�  ��
   ��  1       ��T       ���� $�����  �  �         ����  9 :          "x`� �     �  �  ��
   ��  1       ��T       ���� +�����  �  �         ����  ; <          (h� �     �  ή  ��
   ��  1       ��T       ���� 3�����  �  �         ����  = >          .�p�     @  ��   	   ��  1	       ��T       ���� <U  �  �  �         ����  7 8          ��� � �     �  j�  6+   ��  A        ��U        ���� �����  �  �         ����  9 :          ��� � �     (  �  �C   ��  A       ��U        ���� �����  �  �         ����  ; <          ��� � �     g  ��  n\   ��  A       ��U        ���� �����  �  �         ����  = >          ��� � �     �  V�  
u   ��  A       ��U       ���� �����  �  �         ����  ? @          ��� � �     �  ��  ��   ��  A       ��U       ���� �����  �  �         ����  A B          ��� � �     $  ��  B�   ��  A       ��U       ���� �����  �  �         ����  D E          ��� � �     c  B�  ޾   ��  A       ��U       ���� �����  �  �         ����  F G          ��� � �     �  �  z�   ��  A       ��U       ���� �����  �  �         ����  H I          ��� � �     �  ��  �   ��  A       ��U       ���� &�����  �  �         ����  J K          ��� � �        .�  �	   ��  A	       ��U       ���� /K  �  �  �         ����  ; <          ��� � �     �  ��  �
   ��  B        ��V        ���� �����  �  �         ����  = >          ��� � �        ��   (
   ��  B       ��V        ���� �����  �  �         ����  ? @          ��� � �     H  B�   D
   ��  B       ��V        ���� �����  �  �         ����  A B          ��� � �     �  �  @`
   ��  B       ��V       ���� �����  �  �         ����  C D          ��� � �     �  Ƨ  `|
   ��  B       ��V       ���� �����  �  �         ����  E F          ��� � �        ��  ��
   ��  B       ��V       ���� �����  �  �         ����  H I          ��� � �     h  J�  ��
   ��  B       ��V       ���� $�����  �  �         ����  J K          ��� � �     �  �  ��
   ��  B       ��V       ���� +�����  �  �         ����  L M          ��� �     �  ή  ��
   ��  B       ��V       ���� 3�����  �  �         ����  N O          ��� �     @  ��   	   ��  B	       ��V       ���� <U  �  �  �         ����   5 6          � !�� �     �  j�  6+   ��  R        ��W        ���� �����  �  �         ����   7 8          � '�� �     (  �  �C   ��  R       ��W        ���� �����  �  �         ����   9 :          � -� �     g  ��  n\   ��  R       ��W        ���� �����  �  �         ����   ; <          � 3� �     �  V�  
u   ��  R       ��W       ���� �����  �  �         ����   = >          � 9� �     �  ��  ��   ��  R       ��W       ���� �����  �  �         ����   ? @          � ?� �     $  ��  B�   ��  R       ��W       ���� �����  �  �         ����   B C          � E$� �     c  B�  ޾   ��  R       ��W       ���� �����  �  �         ����   D E          � K,� �     �  �  z�   ��  R       ��W       ���� �����  �  �         ����   F G           Q4� �     �  ��  �   ��  R       ��W       ���� &�����  �  �         ����   H I          W<� �        .�  �	   ��  R	       ��W       ���� /K  �  �  �         ����   9 :          � >"� �     �  ��  �
   ��  S        ��X        ���� �����  �  �         ����   ; <          � E*� �        ��   (
   ��  S       ��X        ���� �����  �  �         ����   = >          � L2� �     H  B�   D
   ��  S       ��X        ���� �����  �  �         ����   ? @          S:� �     �  �  @`
   ��  S       ��X       ���� �����  �  �         ����   A B          ZB� �     �  Ƨ  `|
   ��  S       ��X       ���� �����  �  �         ����   C D          aJ� �        ��  ��
   ��  S       ��X       ���� �����  �  �         ����   F G          hR� �     h  J�  ��
   ��  S       ��X       ���� $�����  �  �         ����   H I          oZ� �     �  �  ��
   ��  S       ��X       ���� +�����  �  �         ����   J K           vb� �     �  ή  ��
   ��  S       ��X       ���� 3�����  �  �         ����   L M          &}j� �     @  ��   	   ��  S	       ��X       ���� <U  �  �  �         ����  D E          �5� � �     �  r�  ��   ��  c        ��Y        ���� �����  �  �         ����  F G          �<� � �     6  �  J�   ��  c       ��Y        ���� �����  �  �         ����  H I          �C� � �     u  ��  ��   ��  c       ��Y        ���� �����  �  �         ����  K L          J� � �     �  ^�  ��   ��  c       ��Y       ���� �����  �  �         ����  M N          Q� � �     �  �  �   ��  c       ��Y       ���� �����  �  �         ����  O P          X� � �     2  ��  �	   ��  c       ��Y       ���� �����  �  �         ����  Q R          _� � �     q  J�  V(	   ��  c       ��Y       ���� �����  �  �         ����  S T          #f� � �     �  �  �@	   ��  c       ��Y       ���� �����  �  �         ����  V W          +m� � �     �  ��  �Y	   ��  c       ��Y       ���� &�����  �  �         ����  X Y          3t� � �     .  6�  *r	   ��  c	       ��Y       ���� /K  �  �  �         ����  I J          [� � �     �  Ƨ  `|
   ��  d        ��Z        ���� �����  �  �         ����  K L          !b� � �        ��  ��
   ��  d       ��Z        ���� �����  �  �         ����  M N          )i� � �     h  J�  ��
   ��  d       ��Z        ���� �����  �  �         ����  P Q          1p� � �     �  �  ��
   ��  d       ��Z       ���� �����  �  �         ����  R S          9w� � �     �  ή  ��
   ��  d       ��Z       ���� �����  �  �         ����  T U          A~� � �     @  ��   	   ��  d       ��Z       ���� �����  �  �         ����  V W          I�� � �     �  R�   %   ��  d       ��Z       ���� $�����  �  �         ����  X Y          Q�� � �     �  �  @A   ��  d       ��Z       ���� +�����  �  �         ����  [ \          Y�� �       ֵ  `]   ��  d       ��Z       ���� 3�����  �  �         ����  ] ^          a�� �     `  ��  �y   ��  d	       ��Z       ���� <U  �  �  �         ����  6 7          � �� �     �  r�  ��   ��  t        ��[        ���� �����  �  �         ����  8 9          � �� �     6  �  J�   ��  t       ��[        ���� �����  �  �         ����  : ;          � %�� �     u  ��  ��   ��  t       ��[        ���� �����  �  �         ����  < =          � +�� �     �  ^�  ��   ��  t       ��[       ���� �����  �  �         ����  > ?          � 1� �     �  �  �   ��  t       ��[       ���� �����  �  �         ����  @ A          � 7� �     2  ��  �	   ��  t       ��[       ���� �����  �  �         ����  C D          � =� �     q  J�  V(	   ��  t       ��[       ���� �����  �  �         ����  E F          � C� �     �  �  �@	   ��  t       ��[       ���� �����  �  �         ����  G H          � I$� �     �  ��  �Y	   ��  t       ��[       ���� &�����  �  �         ����  I J           O,� �     .  6�  *r	   ��  t	       ��[       ���� /K  �  �  �         ����  : ;          � 6� �     �  Ƨ  `|
   ��  u        ��\        ���� �����  �  �         ����  < =          � =� �        ��  ��
   ��  u       ��\        ���� �����  �  �         ����  > ?          � D"� �     h  J�  ��
   ��  u       ��\        ���� �����  �  �         ����  @ A          � K*� �     �  �  ��
   ��  u       ��\       ���� �����  �  �         ����  B C          R2� �     �  ή  ��
   ��  u       ��\       ���� �����  �  �         ����  D E          Y:� �     @  ��   	   ��  u       ��\       ���� �����  �  �         ����  G H          `B� �     �  R�   %   ��  u       ��\       ���� $�����  �  �         ����  I J          gJ� �     �  �  @A   ��  u       ��\       ���� +�����  �  �         ����  K L          nR� �       ֵ  `]   ��  u       ��\       ���� 3�����  �  �         ����  M N           uZ�     `  ��  �y   ��  u	       ��\       ���� <U  �  �  �         ����  5 6          �� �� �     �  r�  ��   ��  �        ��]        ���� �����  �  �         ����  7 8          �� �� �     6  �  J�   ��  �       ��]        ���� �����  �  �         ����  9 :          �� �� �     u  ��  ��   ��  �       ��]        ���� �����  �  �         ����  ; <          �� �� �     �  ^�  ��   ��  �       ��]       ���� �����  �  �         ����  = >          �� �� �     �  �  �   ��  �       ��]       ���� �����  �  �         ����  ? @          �� �� �     2  ��  �	   ��  �       ��]       ���� �����  �  �         ����  B C          �� �� �     q  J�  V(	   ��  �       ��]       ���� �����  �  �         ����  D E          �� �� �     �  �  �@	   ��  �       ��]       ���� �����  �  �         ����  F G          �� �� �     �  ��  �Y	   ��  �       ��]       ���� &�����  �  �         ����  H I          �� �� �     .  6�  *r	   ��  �	       ��]       ���� /K  �  �  �         ����  9 :          �� �� �     �  Ƨ  `|
   ��  �        ��^        ���� �����  �  �         ����  ; <          �� �� �        ��  ��
   ��  �       ��^        ���� �����  �  �         ����  = >          �� �� �     h  J�  ��
   ��  �       ��^        ���� �����  �  �         ����  ? @          �� �� �     �  �  ��
   ��  �       ��^       ���� �����  �  �         ����  A B          �� �� �     �  ή  ��
   ��  �       ��^       ���� �����  �  �         ����  C D          �� �� �     @  ��   	   ��  �       ��^       ���� �����  �  �         ����  F G          �� �� �     �  R�   %   ��  �       ��^       ���� $�����  �  �         ����  H I          �� �� �     �  �  @A   ��  �       ��^       ���� +�����  �  �         ����  J K          �� �� �       ֵ  `]   ��  �       ��^       ���� 3�����  �  �         ����  L M          �� �� �     `  ��  �y   ��  �	       ��^       ���� <U  �  �  �         ����  ( )          � �� �     �  r�  ��   ��  �        ��_        ���� �����  �  �         ����  * +          � "�� �     6  �  J�   ��  �       ��_        ���� �����  �  �         ����  , -          � (� �     u  ��  ��   ��  �       ��_        ���� �����  �  �         ����  . /          � .� �     �  ^�  ��   ��  �       ��_       ���� �����  �  �         ����  0 1          � 4� �     �  �  �   ��  �       ��_       ���� �����  �  �         ����  2 3          � :� �     2  ��  �	   ��  �       ��_       ���� �����  �  �         ����  4 5          � @$� �     q  J�  V(	   ��  �       ��_       ���� �����  �  �         ����  6 7          � F,� �     �  �  �@	   ��  �       ��_       ���� �����  �  �         ����  8 9          � L4� �     �  ��  �Y	   ��  �       ��_       ���� &�����  �  �         ����  : ;          � R<� �     .  6�  *r	   ��  �	       ��_       ���� /K  �  �  �         ����  + ,          � 9"� �     �  Ƨ  `|
   ��  �        ��`        ���� �����  �  �         ����  - .          � @*� �        ��  ��
   ��  �       ��`        ���� �����  �  �         ����  / 0          � G2� �     h  J�  ��
   ��  �       ��`        ���� �����  �  �         ����  1 2          � N:� �     �  �  ��
   ��  �       ��`       ���� �����  �  �         ����  3 4          � UB� �     �  ή  ��
   ��  �       ��`       ���� �����  �  �         ����  5 6          \J� �     @  ��   	   ��  �       ��`       ���� �����  �  �         ����  7 8          cR� �     �  R�   %   ��  �       ��`       ���� $�����  �  �         ����  9 :          jZ� �     �  �  @A   ��  �       ��`       ���� +�����  �  �         ����  ; <          qb� �       ֵ  `]   ��  �       ��`       ���� 3�����  �  �         ����  = >          xj� �     `  ��  �y   ��  �	       ��`       ���� <U  �  �  �         ����  7 8          ��� � �     �  r�  ��   ��  �        ��a        ���� �����  �  �         ����  9 :          ��� � �     6  �  J�   ��  �       ��a        ���� �����  �  �         ����  ; <          ��� � �     u  ��  ��   ��  �       ��a        ���� �����  �  �         ����  = >          ��� � �     �  ^�  ��   ��  �       ��a       ���� �����  �  �         ����  ? @          ��� � �     �  �  �   ��  �       ��a       ���� �����  �  �         ����  A B          ��� � �     2  ��  �	   ��  �       ��a       ���� �����  �  �         ����  D E          ��� � �     q  J�  V(	   ��  �       ��a       ���� �����  �  �         ����  F G          ��� � �     �  �  �@	   ��  �       ��a       ���� �����  �  �         ����  H I          ��� � �     �  ��  �Y	   ��  �       ��a       ���� &�����  �  �         ����  J K          ��� � �     .  6�  *r	   ��  �	       ��a       ���� /K  �  �  �         ����  ; <          ��� � �     �  Ƨ  `|
   ��  �        ��b        ���� �����  �  �         ����  = >          ��� � �        ��  ��
   ��  �       ��b        ���� �����  �  �         ����  ? @          ��� � �     h  J�  ��
   ��  �       ��b        ���� �����  �  �         ����  A B          ��� � �     �  �  ��
   ��  �       ��b       ���� �����  �  �         ����  C D          ��� � �     �  ή  ��
   ��  �       ��b       ���� �����  �  �         ����  E F          ��� � �     @  ��   	   ��  �       ��b       ���� �����  �  �         ����  H I          ��� � �     �  R�   %   ��  �       ��b       ���� $�����  �  �         ����  J K          ��� � �     �  �  @A   ��  �       ��b       ���� +�����  �  �         ����  L M          ��� �       ֵ  `]   ��  �       ��b       ���� 3�����  �  �         ����  N O          ��� �     `  ��  �y   ��  �	       ��b       ���� <U  �  �  �         ����   5 6          � !�� �     �  r�  ��   ��  �        ��c        ���� �����  �  �         ����   7 8          � '�� �     6  �  J�   ��  �       ��c        ���� �����  �  �         ����   9 :          � -�� �     u  ��  ��   ��  �       ��c        ���� �����  �  �         ����   ; <          � 3 � �     �  ^�  ��   ��  �       ��c       ���� �����  �  �         ����   = >          � 9� �     �  �  �   ��  �       ��c       ���� �����  �  �         ����   ? @          � ?� �     2  ��  �	   ��  �       ��c       ���� �����  �  �         ����   B C          � E� �     q  J�  V(	   ��  �       ��c       ���� �����  �  �         ����   D E          � K � �     �  �  �@	   ��  �       ��c       ���� �����  �  �         ����   F G           Q(� �     �  ��  �Y	   ��  �       ��c       ���� &�����  �  �         ����   H I          W0� �     .  6�  *r	   ��  �	       ��c       ���� /K  �  �  �         ����   9 :          � >� �     �  Ƨ  `|
   ��  �        ��d        ���� �����  �  �         ����   ; <          � E� �        ��  ��
   ��  �       ��d        ���� �����  �  �         ����   = >          � L&� �     h  J�  ��
   ��  �       ��d        ���� �����  �  �         ����   ? @          S.� �     �  �  ��
   ��  �       ��d       ���� �����  �  �         ����   A B          Z6� �     �  ή  ��
   ��  �       ��d       ���� �����  �  �         ����   C D          a>� �     @  ��   	   ��  �       ��d       ���� �����  �  �         ����   F G          hF� �     �  R�   %   ��  �       ��d       ���� $�����  �  �         ����   H I          oN� �     �  �  @A   ��  �       ��d       ���� +�����  �  �         ����   J K           vV� �       ֵ  `]   ��  �       ��d       ���� 3�����  �  �         ����   L M          &}^� �     `  ��  �y   ��  �	       ��d       ���� <U  �  �  �         ����  G H          5� � �     �  �  >}   ��  �        ��e        ���� �����  �  �         ����  I J          <� � �     �  ��  ڕ   ��  �       ��e        ���� �����  �  �         ����  K L          "C� � �     9  *�  v�   ��  �       ��e        ���� �����  �  �         ����  N O          *J� � �     x  Ε  �   ��  �       ��e       ���� �����  �  �         ����  P Q          2Q� � �     �  r�  ��   ��  �       ��e       ���� �����  �  �         ����  R S          :X� � �     �  �  J�   ��  �       ��e       ���� �����  �  �         ����  T U          B_� � �     5  ��  �	   ��  �       ��e       ���� �����  �  �         ����  V W          Jf� � �     t  ^�  �)	   ��  �       ��e       ���� �����  �  �         ����  Y Z          Rm� � �     �  �  B	   ��  �       ��e       ���� &�����  �  �         ����  [ \          Zt� � �     �  ��  �Z	   ��  �	       ��e       ���� /K  �  �  �         ����  L M          @[� � �     �  6�  `c
   ��  �        ��f        ���� �����  �  �         ����  N O          Hb� � �     �  ��  �
   ��  �       ��f        ���� �����  �  �         ����  P Q          Pi� � �     (  ��  ��
   ��  �       ��f        ���� �����  �  �         ����  S T          Xp� � �     p  |�  ��
   ��  �       ��f       ���� �����  �  �         ����  U V          `w� � �     �  >�  ��
   ��  �       ��f       ���� �����  �  �         ����  W X          h~� � �         �   �
   ��  �       ��f       ���� �����  �  �         ����  Y Z          p�� � �     H  °      ��  �       ��f       ���� $�����  �  �         ����  [ \          x�� � �     �  ��  @(   ��  �       ��f       ���� +�����  �  �         ����  ^ _          ��� �     �  F�  `D   ��  �       ��f       ���� 3�����  �  �         ����  ` a          ��� �        �  �`   ��  �	       ��f       ���� <U  �  �  �         ����  7 8          � @� �     �  �  >}   ��  �        ��g        ���� �����  �  �         ����  9 :          � F� �     �  ��  ڕ   ��  �       ��g        ���� �����  �  �         ����  ; <          � L� �     9  *�  v�   ��  �       ��g        ���� �����  �  �         ����  = >          R#� �     x  Ε  �   ��  �       ��g       ���� �����  �  �         ����  ? @          X+� �     �  r�  ��   ��  �       ��g       ���� �����  �  �         ����  A B          ^3� �     �  �  J�   ��  �       ��g       ���� �����  �  �         ����  D E          d;� �     5  ��  �	   ��  �       ��g       ���� �����  �  �         ����  F G          jC� �     t  ^�  �)	   ��  �       ��g       ���� �����  �  �         ����  H I           pK� �     �  �  B	   ��  �       ��g       ���� &�����  �  �         ����  J K          &vS� �     �  ��  �Z	   ��  �	       ��g       ���� /K  �  �  �         ����  ; <          ]9� �     �  6�  `c
   ��  �        ��h        ���� �����  �  �         ����  = >          dA� �     �  ��  �
   ��  �       ��h        ���� �����  �  �         ����  ? @          kI� �     (  ��  ��
   ��  �       ��h        ���� �����  �  �         ����  A B          "rQ� �     p  |�  ��
   ��  �       ��h       ���� �����  �  �         ����  C D          (yY� �     �  >�  ��
   ��  �       ��h       ���� �����  �  �         ����  E F          .�a� �         �   �
   ��  �       ��h       ���� �����  �  �         ����  H I          4�i� �     H  °      ��  �       ��h       ���� $�����  �  �         ����  J K          :�q� �     �  ��  @(   ��  �       ��h       ���� +�����  �  �         ����  L M          @�y� �     �  F�  `D   ��  �       ��h       ���� 3�����  �  �         ����  N O          F���        �  �`   ��  �	       ��h       ���� <U  �  �  �         ����  6 7          �� �� �     �  �  >}   ��  �        ��i        ���� �����  �  �         ����  8 9          �� �� �     �  ��  ڕ   ��  �       ��i        ���� �����  �  �         ����  : ;          �� �� �     9  *�  v�   ��  �       ��i        ���� �����  �  �         ����  < =          �� �� �     x  Ε  �   ��  �       ��i       ���� �����  �  �         ����  > ?          �� �� �     �  r�  ��   ��  �       ��i       ���� �����  �  �         ����  @ A          �� �� �     �  �  J�   ��  �       ��i       ���� �����  �  �         ����  C D          �� �� �     5  ��  �	   ��  �       ��i       ���� �����  �  �         ����  E F          �� �� �     t  ^�  �)	   ��  �       ��i       ���� �����  �  �         ����  G H          �� �� �     �  �  B	   ��  �       ��i       ���� &�����  �  �         ����  I J          �� �� �     �  ��  �Z	   ��  �	       ��i       ���� /K  �  �  �         ����  : ;          �� �� �     �  6�  `c
   ��  �        ��j        ���� �����  �  �         ����  < =          �� �� �     �  ��  �
   ��  �       ��j        ���� �����  �  �         ����  > ?          �� �� �     (  ��  ��
   ��  �       ��j        ���� �����  �  �         ����  @ A          �� �� �     p  |�  ��
   ��  �       ��j       ���� �����  �  �         ����  B C          �� �� �     �  >�  ��
   ��  �       ��j       ���� �����  �  �         ����  D E          � � �         �   �
   ��  �       ��j       ���� �����  �  �         ����  G H          � � �     H  °      ��  �       ��j       ���� $�����  �  �         ����  I J          � � �     �  ��  @(   ��  �       ��j       ���� +�����  �  �         ����  K L          � � �     �  F�  `D   ��  �       ��j       ���� 3�����  �  �         ����  M N          &� &� �        �  �`   ��  �	       ��j       ���� <U  �  �  �         ����  ) *          � 7� �     �  �  >}   ��  �        ��k        ���� �����  �  �         ����  + ,          � =� �     �  ��  ڕ   ��  �       ��k        ���� �����  �  �         ����  - .          � C� �     9  *�  v�   ��  �       ��k        ���� �����  �  �         ����  / 0          � I'� �     x  Ε  �   ��  �       ��k       ���� �����  �  �         ����  1 2          � O/� �     �  r�  ��   ��  �       ��k       ���� �����  �  �         ����  3 4          � U7� �     �  �  J�   ��  �       ��k       ���� �����  �  �         ����  5 6          [?� �     5  ��  �	   ��  �       ��k       ���� �����  �  �         ����  7 8          aG� �     t  ^�  �)	   ��  �       ��k       ���� �����  �  �         ����  9 :          gO� �     �  �  B	   ��  �       ��k       ���� &�����  �  �         ����  ; <          mW� �     �  ��  �Z	   ��  �	       ��k       ���� /K  �  �  �         ����  , -          � T=� �     �  6�  `c
   ��  �        ��l        ���� �����  �  �         ����  . /          [E� �     �  ��  �
   ��  �       ��l        ���� �����  �  �         ����  0 1          
bM� �     (  ��  ��
   ��  �       ��l        ���� �����  �  �         ����  2 3          iU� �     p  |�  ��
   ��  �       ��l       ���� �����  �  �         ����  4 5          p]� �     �  >�  ��
   ��  �       ��l       ���� �����  �  �         ����  6 7          we� �         �   �
   ��  �       ��l       ���� �����  �  �         ����  8 9          "~m �     H  °      ��  �       ��l       ���� $�����  �  �         ����  : ;          (�u�     �  ��  @(   ��  �       ��l       ���� +�����  �  �         ����  < =          .�}�     �  F�  `D   ��  �       ��l       ���� 3�����  �  �         ����  > ?          4���        �  �`   ��  �	       ��l       ���� <U  �  �  �         ����  9 :          ��� � �     �  �  >}   ��          ��m        ���� �����  �            ����  ; <          ��� � �     �  ��  ڕ   ��         ��m        ���� �����  �            ����  = >          ��� � �     9  *�  v�   ��         ��m        ���� �����  �            ����  ? @          ��� � �     x  Ε  �   ��         ��m       ���� �����  �            ����  A B          ��� � �     �  r�  ��   ��         ��m       ���� �����  �            ����  C D          ��� � �     �  �  J�   ��         ��m       ���� �����  �            ����  F G          ��� � �     5  ��  �	   ��         ��m       ���� �����  �            ����  H I          ��� � �     t  ^�  �)	   ��         ��m       ���� �����  �            ����  J K          ��� � �     �  �  B	   ��         ��m       ���� &�����  �            ����  L M          ��� � �     �  ��  �Z	   ��  	       ��m       ���� /K  �  �            ����  = >          ��� � �     �  6�  `c
   ��          ��n        ���� �����  �           ����  ? @          ��� � �     �  ��  �
   ��         ��n        ���� �����  �           ����  A B          ��� � �     (  ��  ��
   ��         ��n        ���� �����  �           ����  C D          ��� � �     p  |�  ��
   ��         ��n       ���� �����  �           ����  E F          ��� � �     �  >�  ��
   ��         ��n       ���� �����  �           ����  G H          ��� � �         �   �
   ��         ��n       ���� �����  �           ����  J K          ��� � �     H  °      ��         ��n       ���� $�����  �           ����  L M          ��� � �     �  ��  @(   ��         ��n       ���� +�����  �           ����  N O          �� �     �  F�  `D   ��         ��n       ���� 3�����  �           ����  P Q          �	� �        �  �`   ��  	       ��n       ���� <U  �  �           ����   6 7          � ! � �     �  �  >}   ��          ��o        ���� �����  �           ����   8 9          � '� �     �  ��  ڕ   ��         ��o        ���� �����  �           ����   : ;          � -� �     9  *�  v�   ��         ��o        ���� �����  �           ����   < =          � 3� �     x  Ε  �   ��         ��o       ���� �����  �           ����   > ?          � 9 � �     �  r�  ��   ��         ��o       ���� �����  �           ����   @ A          � ?(� �     �  �  J�   ��         ��o       ���� �����  �           ����   C D          � E0� �     5  ��  �	   ��         ��o       ���� �����  �           ����   E F          � K8� �     t  ^�  �)	   ��         ��o       ���� �����  �           ����   G H           Q@� �     �  �  B	   ��         ��o       ���� &�����  �           ����   I J          WH� �     �  ��  �Z	   ��  	       ��o       ���� /K  �  �           ����   : ;          � >.� �     �  6�  `c
   ��          ��p        ���� �����  �           ����   < =          � E6� �     �  ��  �
   ��         ��p        ���� �����  �           ����   > ?          � L>� �     (  ��  ��
   ��         ��p        ���� �����  �           ����   @ A          SF� �     p  |�  ��
   ��         ��p       ���� �����  �           ����   B C          ZN� �     �  >�  ��
   ��         ��p       ���� �����  �           ����   D E          aV� �         �   �
   ��         ��p       ���� �����  �           ����   G H          h^� �     H  °      ��         ��p       ���� $�����  �           ����   I J          of� �     �  ��  @(   ��         ��p       ���� +�����  �           ����   K L           vn� �     �  F�  `D   ��         ��p       ���� 3�����  �           ����   M N          &}v� �        �  �`   ��  	       ��p       ���� <U  �  �           ����  E F          �5� � �       R�  �e   ��  /        ��q        ���� �����  �           ����  G H           <� � �     �  ��  j~   ��  /       ��q        ���� �����  �           ����  I J          C� � �     �  ��  �   ��  /       ��q        ���� �����  �           ����  L M          J� � �     <  >�  ��   ��  /       ��q       ���� �����  �           ����  N O          Q� � �     {  �  >�   ��  /       ��q       ���� �����  �           ����  P Q           X� � �     �  ��  ��   ��  /       ��q       ���� �����  �           ����  R S          (_� � �     �  *�  v�   ��  /       ��q       ���� �����  �           ����  T U          0f� � �     8  Κ  	   ��  /       ��q       ���� �����  �           ����  W X          8m� � �     w  r�  �*	   ��  /       ��q       ���� &�����  �           ����  Y Z          @t� � �     �  �  JC	   ��  /	       ��q       ���� /K  �  �           ����  J K          &[� � �     X  ��  `J
   ��  0        ��r        ���� �����  �           ����  L M          .b� � �     �  h�  �f
   ��  0       ��r        ���� �����  �           ����  N O          6i� � �     �  *�  ��
   ��  0       ��r        ���� �����  �           ����  Q R          >p� � �     0  �  ��
   ��  0       ��r       ���� �����  �           ����  S T          Fw� � �     x  ��  �
   ��  0       ��r       ���� �����  �           ����  U V          N~� � �     �  p�   �
   ��  0       ��r       ���� �����  �           ����  W X          V�� � �       2�   �
   ��  0       ��r       ���� $�����  �           ����  Y Z          ^�� � �     P  ��  @   ��  0       ��r       ���� +�����  �           ����  \ ]          f�� �     �  ��  `+   ��  0       ��r       ���� 3�����  �           ����  ^ _          n�� �     �  x�  �G   ��  0	       ��r       ���� <U  �  �           ����  6 7          � &�� �       R�  �e   ��  @        ��s        ���� �����  �           ����  8 9          � ,�� �     �  ��  j~   ��  @       ��s        ���� �����  �           ����  : ;          � 2� �     �  ��  �   ��  @       ��s        ���� �����  �           ����  < =          � 8	� �     <  >�  ��   ��  @       ��s       ���� �����  �           ����  > ?          � >� �     {  �  >�   ��  @       ��s       ���� �����  �           ����  @ A          � D� �     �  ��  ��   ��  @       ��s       ���� �����  �           ����  C D          � J!� �     �  *�  v�   ��  @       ��s       ���� �����  �           ����  E F          P)� �     8  Κ  	   ��  @       ��s       ���� �����  �           ����  G H          V1� �     w  r�  �*	   ��  @       ��s       ���� &�����  �           ����  I J          \9� �     �  �  JC	   ��  @	       ��s       ���� /K  �  �           ����  : ;          � C� �     X  ��  `J
   ��  A        ��t        ���� �����  �           ����  < =          � J'� �     �  h�  �f
   ��  A       ��t        ���� �����  �           ����  > ?          Q/� �     �  *�  ��
   ��  A       ��t        ���� �����  �           ����  @ A          	X7� �     0  �  ��
   ��  A       ��t       ���� �����  �           ����  B C          _?� �     x  ��  �
   ��  A       ��t       ���� �����  �           ����  D E          fG� �     �  p�   �
   ��  A       ��t       ���� �����  �           ����  G H          mO� �       2�   �
   ��  A       ��t       ���� $�����  �           ����  I J          !tW� �     P  ��  @   ��  A       ��t       ���� +�����  �           ����  K L          '{_� �     �  ��  `+   ��  A       ��t       ���� 3�����  �           ����  M N          -�g�     �  x�  �G   ��  A	       ��t       ���� <U  �  �           ����  5 6          �� �� �       R�  �e   ��  Q        ��u        ���� �����  �           ����  7 8          �� �� �     �  ��  j~   ��  Q       ��u        ���� �����  �           ����  9 :          �� �� �     �  ��  �   ��  Q       ��u        ���� �����  �           ����  ; <          �� �� �     <  >�  ��   ��  Q       ��u       ���� �����  �           ����  = >          �� �� �     {  �  >�   ��  Q       ��u       ���� �����  �           ����  ? @          �� �� �     �  ��  ��   ��  Q       ��u       ���� �����  �           ����  B C          �� �� �     �  *�  v�   ��  Q       ��u       ���� �����  �           ����  D E          �� �� �     8  Κ  	   ��  Q       ��u       ���� �����  �           ����  F G          �� �� �     w  r�  �*	   ��  Q       ��u       ���� &�����  �           ����  H I          �� �� �     �  �  JC	   ��  Q	       ��u       ���� /K  �  �           ����  9 :          �� �� �     X  ��  `J
   ��  R        ��v        ���� �����  �  	         ����  ; <          �� �� �     �  h�  �f
   ��  R       ��v        ���� �����  �  	         ����  = >          �� �� �     �  *�  ��
   ��  R       ��v        ���� �����  �  	         ����  ? @          �� �� �     0  �  ��
   ��  R       ��v       ���� �����  �  	         ����  A B          �� �� �     x  ��  �
   ��  R       ��v       ���� �����  �  	         ����  C D          �� �� �     �  p�   �
   ��  R       ��v       ���� �����  �  	         ����  F G          �� �� �       2�   �
   ��  R       ��v       ���� $�����  �  	         ����  H I          �� �� �     P  ��  @   ��  R       ��v       ���� +�����  �  	         ����  J K          � � �     �  ��  `+   ��  R       ��v       ���� 3�����  �  	         ����  L M          � � �     �  x�  �G   ��  R	       ��v       ���� <U  �  �  	         ����  ( )          � .� �       R�  �e   ��  b        ��w        ���� �����  �  
         ����  * +          � 4� �     �  ��  j~   ��  b       ��w        ���� �����  �  
         ����  , -          � :� �     �  ��  �   ��  b       ��w        ���� �����  �  
         ����  . /          � @� �     <  >�  ��   ��  b       ��w       ���� �����  �  
         ����  0 1          � F&� �     {  �  >�   ��  b       ��w       ���� �����  �  
         ����  2 3          � L.� �     �  ��  ��   ��  b       ��w       ���� �����  �  
         ����  4 5          � R6� �     �  *�  v�   ��  b       ��w       ���� �����  �  
         ����  6 7          � X>� �     8  Κ  	   ��  b       ��w       ���� �����  �  
         ����  8 9          ^F� �     w  r�  �*	   ��  b       ��w       ���� &�����  �  
         ����  : ;          dN� �     �  �  JC	   ��  b	       ��w       ���� /K  �  �  
         ����  + ,          � K4� �     X  ��  `J
   ��  c        ��x        ���� �����  �           ����  - .          � R<� �     �  h�  �f
   ��  c       ��x        ���� �����  �           ����  / 0          YD� �     �  *�  ��
   ��  c       ��x        ���� �����  �           ����  1 2          `L� �     0  �  ��
   ��  c       ��x       ���� �����  �           ����  3 4          gT� �     x  ��  �
   ��  c       ��x       ���� �����  �           ����  5 6          n\� �     �  p�   �
   ��  c       ��x       ���� �����  �           ����  7 8          ud� �       2�   �
   ��  c       ��x       ���� $�����  �           ����  9 :          |l� �     P  ��  @   ��  c       ��x       ���� +�����  �           ����  ; <          %�t�     �  ��  `+   ��  c       ��x       ���� 3�����  �           ����  = >          +�|	�     �  x�  �G   ��  c	       ��x       ���� <U  �  �           ����  8 9          ��� � �       R�  �e   ��  s        ��y        ���� �����  �           ����  : ;          ��� � �     �  ��  j~   ��  s       ��y        ���� �����  �           ����  < =          ��� � �     �  ��  �   ��  s       ��y        ���� �����  �           ����  > ?          ��� � �     <  >�  ��   ��  s       ��y       ���� �����  �           ����  @ A          ��� � �     {  �  >�   ��  s       ��y       ���� �����  �           ����  B C          ��� � �     �  ��  ��   ��  s       ��y       ���� �����  �           ����  E F          ��� � �     �  *�  v�   ��  s       ��y       ���� �����  �           ����  G H          ��� � �     8  Κ  	   ��  s       ��y       ���� �����  �           ����  I J          ��� � �     w  r�  �*	   ��  s       ��y       ���� &�����  �           ����  K L          ��� � �     �  �  JC	   ��  s	       ��y       ���� /K  �  �           ����  < =          ��� � �     X  ��  `J
   ��  t        ��z        ���� �����  �           ����  > ?          ��� � �     �  h�  �f
   ��  t       ��z        ���� �����  �           ����  @ A          ��� � �     �  *�  ��
   ��  t       ��z        ���� �����  �           ����  B C          ��� � �     0  �  ��
   ��  t       ��z       ���� �����  �           ����  D E          ��� � �     x  ��  �
   ��  t       ��z       ���� �����  �           ����  F G          ��� � �     �  p�   �
   ��  t       ��z       ���� �����  �           ����  I J          ��� � �       2�   �
   ��  t       ��z       ���� $�����  �           ����  K L          ��� � �     P  ��  @   ��  t       ��z       ���� +�����  �           ����  M N          ��� �     �  ��  `+   ��  t       ��z       ���� 3�����  �           ����  O P          ��� �     �  x�  �G   ��  t	       ��z       ���� <U  �  �           ����   5 6          � !�� �       R�  �e   ��  �        ��{        ���� �����  �           ����   7 8          � '�� �     �  ��  j~   ��  �       ��{        ���� �����  �           ����   9 :          � - � �     �  ��  �   ��  �       ��{        ���� �����  �           ����   ; <          � 3� �     <  >�  ��   ��  �       ��{       ���� �����  �           ����   = >          � 9� �     {  �  >�   ��  �       ��{       ���� �����  �           ����   ? @          � ?� �     �  ��  ��   ��  �       ��{       ���� �����  �           ����   B C          � E � �     �  *�  v�   ��  �       ��{       ���� �����  �           ����   D E          � K(� �     8  Κ  	   ��  �       ��{       ���� �����  �           ����   F G           Q0� �     w  r�  �*	   ��  �       ��{       ���� &�����  �           ����   H I          W8� �     �  �  JC	   ��  �	       ��{       ���� /K  �  �           ����   9 :          � >� �     X  ��  `J
   ��  �        ��|        ���� �����  �           ����   ; <          � E&� �     �  h�  �f
   ��  �       ��|        ���� �����  �           ����   = >          � L.� �     �  *�  ��
   ��  �       ��|        ���� �����  �           ����   ? @          S6� �     0  �  ��
   ��  �       ��|       ���� �����  �           ����   A B          Z>� �     x  ��  �
   ��  �       ��|       ���� �����  �           ����   C D          aF� �     �  p�   �
   ��  �       ��|       ���� �����  �           ����   F G          hN� �       2�   �
   ��  �       ��|       ���� $�����  �           ����   H I          oV� �     P  ��  @   ��  �       ��|       ���� +�����  �           ����   J K           v^� �     �  ��  `+   ��  �       ��|       ���� 3�����  �           ����   L M          &}f� �     �  x�  �G   ��  �	       ��|       ���� <U  �  �           ����  F G          
5� � �     3  �  �   ��  �      �   }        ���� �����  �           ����  H I          <� � �     r  ��  ��   ��  �     �   }        ���� �����  �           ����  J K          C� � �     �  J�  V�   ��  �     �   }        ���� �����  �           ����  M N          "J� � �     �  �  ��   ��  �     �   }       ���� �����  �           ����  O P          *Q� � �     /  ��  �	   ��  �     �   }       ���� �����  �           ����  Q R          2X� � �     n  6�  *'	   ��  �     �   }       ���� �����  �           ����  S T          :_� � �     �  ڝ  �?	   ��  �     �   }       ���� �����  �           ����  U V          Bf� � �     �  ~�  bX	   ��  �     �   }       ���� �����  �           ����  X Y          Jm� � �     +  "�  �p	   ��  �     �   }       ���� &�����  �           ����  Z [          Rt� � �     j  Ƣ  ��	   ��  �	     �   }       ���� /K  �  �           ����  K L          8[� � �       V�  `�
   ��  �      �   ~        ���� �����  �           ����  M N          @b� � �     `  �  ��
   ��  �     �   ~        ���� �����  �           ����  O P          Hi� � �     �  ڬ  ��
   ��  �     �   ~        ���� �����  �           ����  R S          Pp� � �     �  ��  ��
   ��  �     �   ~       ���� �����  �           ����  T U          Xw� � �     8  ^�  �   ��  �     �   ~       ���� �����  �           ����  V W          `~� � �     �   �   "   ��  �     �   ~       ���� �����  �           ����  X Y          h�� � �     �  �   >   ��  �     �   ~       ���� $�����  �           ����  Z [          p�� � �       ��  @Z   ��  �     �   ~       ���� +�����  �           ����  ] ^          x�� �     X  f�  `v   ��  �     �   ~       ���� 3�����  �           ����  _ `          ��� �     �  (�  ��   ��  �	     �   ~       ���� <U  �  �           ����  7 8          � 8� �     3  �  �   ��  �      �           ���� �����  �           ����  9 :          � >� �     r  ��  ��   ��  �     �           ���� �����  �           ����  ; <          � D� �     �  J�  V�   ��  �     �           ���� �����  �           ����  = >          � J� �     �  �  ��   ��  �     �          ���� �����  �           ����  ? @           P#� �     /  ��  �	   ��  �     �          ���� �����  �           ����  A B          V+� �     n  6�  *'	   ��  �     �          ���� �����  �           ����  D E          \3� �     �  ڝ  �?	   ��  �     �          ���� �����  �           ����  F G          b;� �     �  ~�  bX	   ��  �     �          ���� �����  �           ����  H I          hC� �     +  "�  �p	   ��  �     �          ���� &�����  �           ����  J K          nK� �     j  Ƣ  ��	   ��  �	     �          ���� /K  �  �           ����  ; <          U1� �       V�  `�
   ��  �      �   �        ���� �����  �           ����  = >          \9� �     `  �  ��
   ��  �     �   �        ���� �����  �           ����  ? @          cA� �     �  ڬ  ��
   ��  �     �   �        ���� �����  �           ����  A B          jI� �     �  ��  ��
   ��  �     �   �       ���� �����  �           ����  C D           qQ� �     8  ^�  �   ��  �     �   �       ���� �����  �           ����  E F          &xY� �     �   �   "   ��  �     �   �       ���� �����  �           ����  H I          ,a� �     �  �   >   ��  �     �   �       ���� $�����  �           ����  J K          2�i� �       ��  @Z   ��  �     �   �       ���� +�����  �           ����  L M          8�q� �     X  f�  `v   ��  �     �   �       ���� 3�����  �           ����  N O          >�y�     �  (�  ��   ��  �	     �   �       ���� <U  �  �           ����  6 7          �� �� �     3  �  �   ��  �      �   �        ���� �����  �           ����  8 9          �� �� �     r  ��  ��   ��  �     �   �        ���� �����  �           ����  : ;          �� �� �     �  J�  V�   ��  �     �   �        ���� �����  �           ����  < =          �� �� �     �  �  ��   ��  �     �   �       ���� �����  �           ����  > ?          �� �� �     /  ��  �	   ��  �     �   �       ���� �����  �           ����  @ A          �� �� �     n  6�  *'	   ��  �     �   �       ���� �����  �           ����  C D          �� �� �     �  ڝ  �?	   ��  �     �   �       ���� �����  �           ����  E F          �� �� �     �  ~�  bX	   ��  �     �   �       ���� �����  �           ����  G H          �� �� �     +  "�  �p	   ��  �     �   �       ���� &�����  �           ����  I J          �� �� �     j  Ƣ  ��	   ��  �	     �   �       ���� /K  �  �           ����  : ;          �� �� �       V�  `�
   ��  �      �   �        ���� �����  �           ����  < =          �� �� �     `  �  ��
   ��  �     �   �        ���� �����  �           ����  > ?          �� �� �     �  ڬ  ��
   ��  �     �   �        ���� �����  �           ����  @ A          �� �� �     �  ��  ��
   ��  �     �   �       ���� �����  �           ����  B C          �� �� �     8  ^�  �   ��  �     �   �       ���� �����  �           ����  D E          �� �� �     �   �   "   ��  �     �   �       ���� �����  �           ����  G H          � � �     �  �   >   ��  �     �   �       ���� $�����  �           ����  I J          � � �       ��  @Z   ��  �     �   �       ���� +�����  �           ����  K L          � � �     X  f�  `v   ��  �     �   �       ���� 3�����  �           ����  M N          � � �     �  (�  ��   ��  �	     �   �       ���� <U  �  �           ����  * +          � �� �     3  �  �   ��  �      �   �        ���� �����  �           ����  , -          � !�� �     r  ��  ��   ��  �     �   �        ���� �����  �           ����  . /          � '�� �     �  J�  V�   ��  �     �   �        ���� �����  �           ����  0 1          � -� �     �  �  ��   ��  �     �   �       ���� �����  �           ����  2 3          � 3� �     /  ��  �	   ��  �     �   �       ���� �����  �           ����  4 5          � 9� �     n  6�  *'	   ��  �     �   �       ���� �����  �           ����  6 7          � ?� �     �  ڝ  �?	   ��  �     �   �       ���� �����  �           ����  8 9          � E&� �     �  ~�  bX	   ��  �     �   �       ���� �����  �           ����  : ;          � K.� �     +  "�  �p	   ��  �     �   �       ���� &�����  �           ����  < =          Q6� �     j  Ƣ  ��	   ��  �	     �   �       ���� /K  �  �           ����  - .          � 8� �       V�  `�
   ��  �      �   �        ���� �����  �           ����  / 0          � ?$� �     `  �  ��
   ��  �     �   �        ���� �����  �           ����  1 2          � F,� �     �  ڬ  ��
   ��  �     �   �        ���� �����  �           ����  3 4          � M4� �     �  ��  ��
   ��  �     �   �       ���� �����  �           ����  5 6          T<� �     8  ^�  �   ��  �     �   �       ���� �����  �           ����  7 8          
[D� �     �   �   "   ��  �     �   �       ���� �����  �           ����  9 :          bL� �     �  �   >   ��  �     �   �       ���� $�����  �           ����  ; <          iT� �       ��  @Z   ��  �     �   �       ���� +�����  �           ����  = >          p\� �     X  f�  `v   ��  �     �   �       ���� 3�����  �           ����  ? @          "wd �     �  (�  ��   ��  �	     �   �       ���� <U  �  �           ����   6 7          � !�� �     3  �  �   ��  �      �   �        ���� �����  �           ����   8 9          � '� �     r  ��  ��   ��  �     �   �        ���� �����  �           ����   : ;          � -� �     �  J�  V�   ��  �     �   �        ���� �����  �           ����   < =          � 3� �     �  �  ��   ��  �     �   �       ���� �����  �           ����   > ?          � 9� �     /  ��  �	   ��  �     �   �       ���� �����  �           ����   @ A          � ?$� �     n  6�  *'	   ��  �     �   �       ���� �����  �           ����   C D          � E,� �     �  ڝ  �?	   ��  �     �   �       ���� �����  �           ����   E F          � K4� �     �  ~�  bX	   ��  �     �   �       ���� �����  �           ����   G H           Q<� �     +  "�  �p	   ��  �     �   �       ���� &�����  �           ����   I J          WD� �     j  Ƣ  ��	   ��  �	     �   �       ���� /K  �  �           ����   : ;          � >*� �       V�  `�
   ��  �      �   �        ���� �����  �           ����   < =          � E2� �     `  �  ��
   ��  �     �   �        ���� �����  �           ����   > ?          � L:� �     �  ڬ  ��
   ��  �     �   �        ���� �����  �           ����   @ A          SB� �     �  ��  ��
   ��  �     �   �       ���� �����  �           ����   B C          ZJ� �     8  ^�  �   ��  �     �   �       ���� �����  �           ����   D E          aR� �     �   �   "   ��  �     �   �       ���� �����  �           ����   G H          hZ� �     �  �   >   ��  �     �   �       ���� $�����  �           ����   I J          ob� �       ��  @Z   ��  �     �   �       ���� +�����  �           ����   K L           vj� �     X  f�  `v   ��  �     �   �       ���� 3�����  �           ����   M N          &}r� �     �  (�  ��   ��  �	     �   �       ���� <U  �  �           % ��  G H           5� � �     ������  ��       �       �    �        ���� �����  �           % ��  I J           <� � �     ����6�  *�       �      �    �        ���� �����  �           % ��  K L           'C� � �     ����ژ  ��       �      �    �        ���� �����  �           & ��  N O           /J� � �     ����~�  b	       �      �    �        ���� �����  �           & ��  P Q           7Q� � �     ����"�  �%	       �      �    �        ���� �����  �           & ��  R S           ?X� � �     ����Ɲ  �>	       �      �    �        ���� �����  �           ' ��  T U           G_� � �     ����j�  6W	       �      �    �        ���� �����  �           ' ��  V W           Of� � �     �����  �o	       �      �    �        ���� �����  �           ' ��  Y Z           Wm� � �     ������  n�	       �      �    �        ���� &�����  �           ( ��  [ \           _t� � �     ����V�  
�	       � 	     �    �        ���� /�����  �           ) ��  L M           E[� � �     �����  `�
       �       �    �        ���� �����  �           ) ��  N O           Mb� � �     ������  ��
       �      �    �        ���� �����  �           ) ��  P Q           Ui� � �     ����j�  ��
       �      �    �        ���� �����  �           * ��  S T           ]p� � �     ����,�  �       �      �    �        ���� �����  �           * ��  U V           ew� � �     �����  �       �      �    �        ���� �����  �           * ��  W X           m~� � �     ������   ;       �      �    �        ���� �����  �           + ��  Y Z           u�� � �     ����r�   W       �      �    �        ���� $�����  �           + ��  [ \           }�� � �     ����4�  @s       �      �    �        ���� +�����  �           + ��  ^ _           ��� �     ������  `�       �      �    �        ���� 3�����  �           , ��  ` a           ��� �     ������  ��       � 	     �    �        ���� <�����  �           % ��  7 8           � E� �     ������  ��       �       �    �        ���� �����  �           % ��  9 :           � K� �     ����6�  *�       �      �    �        ���� �����  �           % ��  ; <           Q � �     ����ژ  ��       �      �    �        ���� �����  �           & ��  = >           W(� �     ����~�  b	       �      �    �        ���� �����  �           & ��  ? @           ]0� �     ����"�  �%	       �      �    �        ���� �����  �           & ��  A B           c8� �     ����Ɲ  �>	       �      �    �        ���� �����  �           ' ��  D E           i@� �     ����j�  6W	       �      �    �        ���� �����  �           ' ��  F G           oH� �     �����  �o	       �      �    �        ���� �����  �           ' ��  H I           %uP� �     ������  n�	       �      �    �        ���� &�����  �           ( ��  J K           +{X� �     ����V�  
�	       � 	     �    �        ���� /�����  �           ) ��  ; <           b>� �     �����  `�
       �       �    �        ���� �����  �           ) ��  = >           iF� �     ������  ��
       �      �    �        ���� �����  �           ) ��  ? @           !pN� �     ����j�  ��
       �      �    �        ���� �����  �           * ��  A B           'wV� �     ����,�  �       �      �    �        ���� �����  �           * ��  C D           -~^� �     �����  �       �      �    �        ���� �����  �           * ��  E F           3�f� �     ������   ;       �      �    �        ���� �����  �           + ��  H I           9�n� �     ����r�   W       �      �    �        ���� $�����  �           + ��  J K           ?�v� �     ����4�  @s       �      �    �        ���� +�����  �           + ��  L M           E�~� �     ������  `�       �      �    �        ���� 3�����  �           , ��  N O           K���     ������  ��       � 	     �    �        ���� <�����  �           % ��  6 7           �� �� �     ������  ��       �       �    �        ���� �����  �           % ��  8 9           �� �� �     ����6�  *�       �      �    �        ���� �����  �           % ��  : ;           �� �� �     ����ژ  ��       �      �    �        ���� �����  �           & ��  < =           �� �� �     ����~�  b	       �      �    �        ���� �����  �           & ��  > ?           �� �� �     ����"�  �%	       �      �    �        ���� �����  �           & ��  @ A           �� �� �     ����Ɲ  �>	       �      �    �        ���� �����  �           ' ��  C D           �� �� �     ����j�  6W	       �      �    �        ���� �����  �           ' ��  E F           �� �� �     �����  �o	       �      �    �        ���� �����  �           ' ��  G H           �� �� �     ������  n�	       �      �    �        ���� &�����  �           ( ��  I J           �� �� �     ����V�  
�	       � 	     �    �        ���� /�����  �           ) ��  : ;           �� �� �     �����  `�
       �       �    �        ���� �����  �           ) ��  < =           �� �� �     ������  ��
       �      �    �        ���� �����  �           ) ��  > ?           �� �� �     ����j�  ��
       �      �    �        ���� �����  �           * ��  @ A           �� �� �     ����,�  �       �      �    �        ���� �����  �           * ��  B C           � � �     �����  �       �      �    �        ���� �����  �           * ��  D E           � � �     ������   ;       �      �    �        ���� �����  �           + ��  G H           � � �     ����r�   W       �      �    �        ���� $�����  �           + ��  I J           � � �     ����4�  @s       �      �    �        ���� +�����  �           + ��  K L           #� #� �     ������  `�       �      �    �        ���� 3�����  �           , ��  M N           +� +� �     ������  ��       � 	     �    �        ���� <�����  �           % ��  ) *           � 0� �     ������  ��       �       �    �        ���� �����  �            % ��  + ,           � 6� �     ����6�  *�       �      �    �        ���� �����  �            % ��  - .           � <� �     ����ژ  ��       �      �    �        ���� �����  �            & ��  / 0           � B� �     ����~�  b	       �      �    �        ���� �����  �            & ��  1 2           � H#� �     ����"�  �%	       �      �    �        ���� �����  �            & ��  3 4           � N+� �     ����Ɲ  �>	       �      �    �        ���� �����  �            ' ��  5 6           T3� �     ����j�  6W	       �      �    �        ���� �����  �            ' ��  7 8           	Z;� �     �����  �o	       �      �    �        ���� �����  �            ' ��  9 :           `C� �     ������  n�	       �      �    �        ���� &�����  �            ( ��  ; <           fK� �     ����V�  
�	       � 	     �    �        ���� /�����  �            ) ��  , -           � M1� �     �����  `�
       �       �    �        ���� �����  �  !         ) ��  . /           T9� �     ������  ��
       �      �    �        ���� �����  �  !         ) ��  0 1           [A� �     ����j�  ��
       �      �    �        ���� �����  �  !         * ��  2 3           bI� �     ����,�  �       �      �    �        ���� �����  �  !         * ��  4 5           iQ� �     �����  �       �      �    �        ���� �����  �  !         * ��  6 7           pY� �     ������   ;       �      �    �        ���� �����  �  !         + ��  8 9           #wa�     ����r�   W       �      �    �        ���� $�����  �  !         + ��  : ;           )~i
�     ����4�  @s       �      �    �        ���� +�����  �  !         + ��  < =           /�q�     ������  `�       �      �    �        ���� 3�����  �  !         , ��  > ?           5�y�     ������  ��       � 	     �    �        ���� <�����  �  !         % ��  8 9           ��� � �     ������  ��             �     �        ���� �����  �  "         % ��  : ;           ��� � �     ����6�  *�            �     �        ���� �����  �  "         % ��  < =           ��� � �     ����ژ  ��            �     �        ���� �����  �  "         & ��  > ?           ��� � �     ����~�  b	            �     �        ���� �����  �  "         & ��  @ A           ��� � �     ����"�  �%	            �     �        ���� �����  �  "         & ��  B C           ��� � �     ����Ɲ  �>	            �     �        ���� �����  �  "         ' ��  E F           ��� � �     ����j�  6W	            �     �        ���� �����  �  "         ' ��  G H           ��� � �     �����  �o	            �     �        ���� �����  �  "         ' ��  I J           ��� � �     ������  n�	            �     �        ���� &�����  �  "         ( ��  K L           ��� � �     ����V�  
�	       	     �     �        ���� /�����  �  "         ) ��  < =           ��� � �     �����  `�
             �     �        ���� �����  �  #         ) ��  > ?           ��� � �     ������  ��
            �     �        ���� �����  �  #         ) ��  @ A           ��� � �     ����j�  ��
            �     �        ���� �����  �  #         * ��  B C           ��� � �     ����,�  �            �     �        ���� �����  �  #         * ��  D E           ��� � �     �����  �            �     �        ���� �����  �  #         * ��  F G           ��� � �     ������   ;            �     �        ���� �����  �  #         + ��  I J           ��� � �     ����r�   W            �     �        ���� $�����  �  #         + ��  K L           ��� � �     ����4�  @s            �     �        ���� +�����  �  #         + ��  M N           �� �     ������  `�            �     �        ���� 3�����  �  #         , ��  O P           �
� �     ������  ��       	     �     �        ���� <�����  �  #         % ��   6 7           � !� �     ������  ��             � !   �        ���� �����  �  $         % ��   8 9           � '� �     ����6�  *�            � !   �        ���� �����  �  $         % ��   : ;           � -� �     ����ژ  ��            � !   �        ���� �����  �  $         & ��   < =           � 3'� �     ����~�  b	            � !   �        ���� �����  �  $         & ��   > ?           � 9/� �     ����"�  �%	            � !   �        ���� �����  �  $         & ��   @ A           � ?7� �     ����Ɲ  �>	            � !   �        ���� �����  �  $         ' ��   C D           � E?� �     ����j�  6W	            � !   �        ���� �����  �  $         ' ��   E F           � KG� �     �����  �o	            � !   �        ���� �����  �  $         ' ��   G H            QO� �     ������  n�	            � !   �        ���� &�����  �  $         ( ��   I J           WW� �     ����V�  
�	       	     � !   �        ���� /�����  �  $         ) ��   : ;           � >=� �     �����  `�
             � !   �        ���� �����  �  %         ) ��   < =           � EE� �     ������  ��
            � !   �        ���� �����  �  %         ) ��   > ?           � LM� �     ����j�  ��
            � !   �        ���� �����  �  %         * ��   @ A           SU� �     ����,�  �            � !   �        ���� �����  �  %         * ��   B C           Z]� �     �����  �            � !   �        ���� �����  �  %         * ��   D E           ae� �     ������   ;            � !   �        ���� �����  �  %         + ��   G H           hm� �     ����r�   W            � !   �        ���� $�����  �  %         + ��   I J           ou� �     ����4�  @s            � !   �        ���� +�����  �  %         + ��   K L            v}� �     ������  `�            � !   �        ���� 3�����  �  %         , ��   M N           &}�� �     ������  ��       	     � !   �        ���� <�����  �  %         ����	  D E           �5� � �     ������  n�   ��  �      �� ���        ���� �����  �  &         ����	  F G           �<� � �     ����V�  
	   ��  �     �� ���        ���� �����  �  &         ����	  H I           C� � �     ������  �#	   ��  �     �� ���        ���� �����  �  &         ����	  K L           J� � �     ������  B<	   ��  �     �� ���       ���� �����  �  &         ����	  M N           Q� � �     ����B�  �T	   ��  �     �� ���       ���� �����  �  &         ����	  O P           X� � �     �����  zm	   ��  �     �� ���       ���� �����  �  &         ����	  Q R           #_� � �     ������  �	   ��  �     �� ���       ���� �����  �  &         ����	  S T           +f� � �     ����.�  ��	   ��  �     �� ���       ���� �����  �  &         ����	  V W           3m� � �     ����ҥ  N�	   ��  �     �� ���       ���� &�����  �  &         ����	  X Y           ;t� � �     ����v�  ��	   ��  �	     �� ���       ���� /�����  �  &         ����	  I J           ![� � �     �����  `�
   ��  �      �� ���        ���� �����  �  '         ����	  K L           )b� � �     ����ȯ  ��
   ��  �     �� ���        ���� �����  �  '         ����	  M N           1i� � �     ������  �   ��  �     �� ���        ���� �����  �  '         ����	  P Q           9p� � �     ����L�  �4   ��  �     �� ���       ���� �����  �  '         ����	  R S           Aw� � �     �����  �P   ��  �     �� ���       ���� �����  �  '         ����	  T U           I~� � �     ����ж   m   ��  �     �� ���       ���� �����  �  '         ����	  V W           Q�� � �     ������   �   ��  �     �� ���       ���� $�����  �  '         ����	  X Y           Y�� � �     ����T�  @�   ��  �     �� ���       ���� +�����  �  '         ����	  [ \           a�� �     �����  `�   ��  �     �� ���       ���� 3�����  �  '         ����	  ] ^           i�� �     ����ؽ  ��   ��  �	     �� ���       ���� <�����  �  '         ����	  6 7           � !�� �     ������  n�   ��  �      �� ���        ���� �����  �  (         ����	  8 9           � '�� �     ����V�  
	   ��  �     �� ���        ���� �����  �  (         ����	  : ;           � -�� �     ������  �#	   ��  �     �� ���        ���� �����  �  (         ����	  < =           � 3� �     ������  B<	   ��  �     �� ���       ���� �����  �  (         ����	  > ?           � 9� �     ����B�  �T	   ��  �     �� ���       ���� �����  �  (         ����	  @ A           � ?� �     �����  zm	   ��  �     �� ���       ���� �����  �  (         ����	  C D           � E� �     ������  �	   ��  �     �� ���       ���� �����  �  (         ����	  E F           � K$� �     ����.�  ��	   ��  �     �� ���       ���� �����  �  (         ����	  G H           Q,� �     ����ҥ  N�	   ��  �     �� ���       ���� &�����  �  (         ����	  I J           W4� �     ����v�  ��	   ��  �	     �� ���       ���� /�����  �  (         ����	  : ;           � >� �     �����  `�
   ��  �      �� ���        ���� �����  �  )         ����	  < =           � E"� �     ����ȯ  ��
   ��  �     �� ���        ���� �����  �  )         ����	  > ?           � L*� �     ������  �   ��  �     �� ���        ���� �����  �  )         ����	  @ A           S2� �     ����L�  �4   ��  �     �� ���       ���� �����  �  )         ����	  B C           
Z:� �     �����  �P   ��  �     �� ���       ���� �����  �  )         ����	  D E           aB� �     ����ж   m   ��  �     �� ���       ���� �����  �  )         ����	  G H           hJ� �     ������   �   ��  �     �� ���       ���� $�����  �  )         ����	  I J           oR� �     ����T�  @�   ��  �     �� ���       ���� +�����  �  )         ����	  K L           "vZ� �     �����  `�   ��  �     �� ���       ���� 3�����  �  )         ����	  M N           (}b�     ����ؽ  ��   ��  �	     �� ���       ���� <�����  �  )         ����	  5 6           �� �� �     ������  n�   ��        �� ���        ���� �����  �  *         ����	  7 8           �� �� �     ����V�  
	   ��       �� ���        ���� �����  �  *         ����	  9 :           �� �� �     ������  �#	   ��       �� ���        ���� �����  �  *         ����	  ; <           �� �� �     ������  B<	   ��       �� ���       ���� �����  �  *         ����	  = >           �� �� �     ����B�  �T	   ��       �� ���       ���� �����  �  *         ����	  ? @           �� �� �     �����  zm	   ��       �� ���       ���� �����  �  *         ����	  B C           �� �� �     ������  �	   ��       �� ���       ���� �����  �  *         ����	  D E           �� �� �     ����.�  ��	   ��       �� ���       ���� �����  �  *         ����	  F G           �� �� �     ����ҥ  N�	   ��       �� ���       ���� &�����  �  *         ����	  H I           �� �� �     ����v�  ��	   ��  	     �� ���       ���� /�����  �  *         ����	  9 :           �� �� �     �����  `�
   ��  	      �� ���        ���� �����  �  +         ����	  ; <           �� �� �     ����ȯ  ��
   ��  	     �� ���        ���� �����  �  +         ����	  = >           �� �� �     ������  �   ��  	     �� ���        ���� �����  �  +         ����	  ? @           �� �� �     ����L�  �4   ��  	     �� ���       ���� �����  �  +         ����	  A B           �� �� �     �����  �P   ��  	     �� ���       ���� �����  �  +         ����	  C D           �� �� �     ����ж   m   ��  	     �� ���       ���� �����  �  +         ����	  F G           �� �� �     ������   �   ��  	     �� ���       ���� $�����  �  +         ����	  H I           �� �� �     ����T�  @�   ��  	     �� ���       ���� +�����  �  +         ����	  J K           �� �� �     �����  `�   ��  	     �� ���       ���� 3�����  �  +         ����	  L M           � � �     ����ؽ  ��   ��  		     �� ���       ���� <�����  �  +         ����	  ) *           � �� �     ������  n�   ��        �� ���        ���� �����  �  ,         ����	  + ,           � �� �     ����V�  
	   ��       �� ���        ���� �����  �  ,         ����	  - .           � $�� �     ������  �#	   ��       �� ���        ���� �����  �  ,         ����	  / 0           � *� �     ������  B<	   ��       �� ���       ���� �����  �  ,         ����	  1 2           � 0� �     ����B�  �T	   ��       �� ���       ���� �����  �  ,         ����	  3 4           � 6� �     �����  zm	   ��       �� ���       ���� �����  �  ,         ����	  5 6           � <� �     ������  �	   ��       �� ���       ���� �����  �  ,         ����	  7 8           � B#� �     ����.�  ��	   ��       �� ���       ���� �����  �  ,         ����	  9 :           � H+� �     ����ҥ  N�	   ��       �� ���       ���� &�����  �  ,         ����	  ; <           N3� �     ����v�  ��	   ��  	     �� ���       ���� /�����  �  ,         ����	  , -           � 5� �     �����  `�
   ��        �� ���        ���� �����  �  -         ����	  . /           � <!� �     ����ȯ  ��
   ��       �� ���        ���� �����  �  -         ����	  0 1           � C)� �     ������  �   ��       �� ���        ���� �����  �  -         ����	  2 3           J1� �     ����L�  �4   ��       �� ���       ���� �����  �  -         ����	  4 5           Q9� �     �����  �P   ��       �� ���       ���� �����  �  -         ����	  6 7           XA� �     ����ж   m   ��       �� ���       ���� �����  �  -         ����	  8 9           _I� �     ������   �   ��       �� ���       ���� $�����  �  -         ����	  : ;           fQ� �     ����T�  @�   ��       �� ���       ���� +�����  �  -         ����	  < =           mY� �     �����  `�   ��       �� ���       ���� 3�����  �  -         ����	  > ?           %ta �     ����ؽ  ��   ��  	     �� ���       ���� <�����  �  -         ����	  7 8           ��� � �     ������  n�   ��  &      ��  ���        ���� �����  �  .         ����	  9 :           ��� � �     ����V�  
	   ��  &     ��  ���        ���� �����  �  .         ����	  ; <           ��� � �     ������  �#	   ��  &     ��  ���        ���� �����  �  .         ����	  = >           ��� � �     ������  B<	   ��  &     ��  ���       ���� �����  �  .         ����	  ? @           ��� � �     ����B�  �T	   ��  &     ��  ���       ���� �����  �  .         ����	  A B           ��� � �     �����  zm	   ��  &     ��  ���       ���� �����  �  .         ����	  D E           ��� � �     ������  �	   ��  &     ��  ���       ���� �����  �  .         ����	  F G           ��� � �     ����.�  ��	   ��  &     ��  ���       ���� �����  �  .         ����	  H I           ��� � �     ����ҥ  N�	   ��  &     ��  ���       ���� &�����  �  .         ����	  J K           ��� � �     ����v�  ��	   ��  &	     ��  ���       ���� /�����  �  .         ����	  ; <           ��� � �     �����  `�
   ��  '      ��  ���        ���� �����  �  /         ����	  = >           ��� � �     ����ȯ  ��
   ��  '     ��  ���        ���� �����  �  /         ����	  ? @           ��� � �     ������  �   ��  '     ��  ���        ���� �����  �  /         ����	  A B           ��� � �     ����L�  �4   ��  '     ��  ���       ���� �����  �  /         ����	  C D           ��� � �     �����  �P   ��  '     ��  ���       ���� �����  �  /         ����	  E F           ��� � �     ����ж   m   ��  '     ��  ���       ���� �����  �  /         ����	  H I           ��� � �     ������   �   ��  '     ��  ���       ���� $�����  �  /         ����	  J K           ��� � �     ����T�  @�   ��  '     ��  ���       ���� +�����  �  /         ����	  L M           ��� �     �����  `�   ��  '     ��  ���       ���� 3�����  �  /         ����	  N O           ��� �     ����ؽ  ��   ��  '	     ��  ���       ���� <�����  �  /         ����	   5 6           � !�� �     ������  n�   ��  5      ��! ���        ���� �����  �  0         ����	   7 8           � '�� �     ����V�  
	   ��  5     ��! ���        ���� �����  �  0         ����	   9 :           � -�� �     ������  �#	   ��  5     ��! ���        ���� �����  �  0         ����	   ; <           � 3� �     ������  B<	   ��  5     ��! ���       ���� �����  �  0         ����	   = >           � 9� �     ����B�  �T	   ��  5     ��! ���       ���� �����  �  0         ����	   ? @           � ?� �     �����  zm	   ��  5     ��! ���       ���� �����  �  0         ����	   B C           � E� �     ������  �	   ��  5     ��! ���       ���� �����  �  0         ����	   D E           � K&� �     ����.�  ��	   ��  5     ��! ���       ���� �����  �  0         ����	   F G            Q.� �     ����ҥ  N�	   ��  5     ��! ���       ���� &�����  �  0         ����	   H I           W6� �     ����v�  ��	   ��  5	     ��! ���       ���� /�����  �  0         ����	   9 :           � >� �     �����  `�
   ��  6      ��! ���        ���� �����  �  1         ����	   ; <           � E$� �     ����ȯ  ��
   ��  6     ��! ���        ���� �����  �  1         ����	   = >           � L,� �     ������  �   ��  6     ��! ���        ���� �����  �  1         ����	   ? @           S4� �     ����L�  �4   ��  6     ��! ���       ���� �����  �  1         ����	   A B           Z<� �     �����  �P   ��  6     ��! ���       ���� �����  �  1         ����	   C D           aD� �     ����ж   m   ��  6     ��! ���       ���� �����  �  1         ����	   F G           hL� �     ������   �   ��  6     ��! ���       ���� $�����  �  1         ����	   H I           oT� �     ����T�  @�   ��  6     ��! ���       ���� +�����  �  1         ����	   J K            v\� �     �����  `�   ��  6     ��! ���       ���� 3�����  �  1         ����	   L M           &}d� �     ����ؽ  ��   ��  6	     ��! ���       ���� <�����  �  1         ����
  E F            5� � �     ����"�  ��   ��  D      �� ���        ���� �����  �  2         ����
  G H           <� � �     ����Ƙ  ��   ��  D     �� ���        ���� �����  �  2         ����
  I J           C� � �     ����j�  6	   ��  D     �� ���        ���� �����  �  2         ����
  L M           J� � �     �����  �$	   ��  D     �� ���       ���� �����  �  2         ����
  N O            Q� � �     ������  n=	   ��  D     �� ���       ���� �����  �  2         ����
  P Q           (X� � �     ����V�  
V	   ��  D     �� ���       ���� �����  �  2         ����
  R S           0_� � �     ������  �n	   ��  D     �� ���       ���� �����  �  2         ����
  T U           8f� � �     ������  B�	   ��  D     �� ���       ���� �����  �  2         ����
  W X           @m� � �     ����B�  ޟ	   ��  D     �� ���       ���� &�����  �  2         ����
  Y Z           Ht� � �     �����  z�	   ��  D	     �� ���       ���� /�����  �  2         ����
  J K           .[� � �     ����v�  `�
   ��  E      �� ���        ���� �����  �  3         ����
  L M           6b� � �     ����8�  ��
   ��  E     �� ���        ���� �����  �  3         ����
  N O           >i� � �     ������  ��
   ��  E     �� ���        ���� �����  �  3         ����
  Q R           Fp� � �     ������  �   ��  E     �� ���       ���� �����  �  3         ����
  S T           Nw� � �     ����~�  �7   ��  E     �� ���       ���� �����  �  3         ����
  U V           V~� � �     ����@�   T   ��  E     �� ���       ���� �����  �  3         ����
  W X           ^�� � �     �����   p   ��  E     �� ���       ���� $�����  �  3         ����
  Y Z           f�� � �     ����ĸ  @�   ��  E     �� ���       ���� +�����  �  3         ����
  \ ]           n�� �     ������  `�   ��  E     �� ���       ���� 3�����  �  3         ����
  ^ _           v�� �     ����H�  ��   ��  E	     �� ���       ���� <�����  �  3         ����
  6 7           � .�� �     ����"�  ��   ��  S      �� ���        ���� �����  �  4         ����
  8 9           � 4� �     ����Ƙ  ��   ��  S     �� ���        ���� �����  �  4         ����
  : ;           � :	� �     ����j�  6	   ��  S     �� ���        ���� �����  �  4         ����
  < =           � @� �     �����  �$	   ��  S     �� ���       ���� �����  �  4         ����
  > ?           � F� �     ������  n=	   ��  S     �� ���       ���� �����  �  4         ����
  @ A           � L!� �     ����V�  
V	   ��  S     �� ���       ���� �����  �  4         ����
  C D           R)� �     ������  �n	   ��  S     �� ���       ���� �����  �  4         ����
  E F           	X1� �     ������  B�	   ��  S     �� ���       ���� �����  �  4         ����
  G H           ^9� �     ����B�  ޟ	   ��  S     �� ���       ���� &�����  �  4         ����
  I J           dA� �     �����  z�	   ��  S	     �� ���       ���� /�����  �  4         ����
  : ;           � K'� �     ����v�  `�
   ��  T      �� ���        ���� �����  �  5         ����
  < =           R/� �     ����8�  ��
   ��  T     �� ���        ���� �����  �  5         ����
  > ?           Y7� �     ������  ��
   ��  T     �� ���        ���� �����  �  5         ����
  @ A           `?� �     ������  �   ��  T     �� ���       ���� �����  �  5         ����
  B C           gG� �     ����~�  �7   ��  T     �� ���       ���� �����  �  5         ����
  D E           nO� �     ����@�   T   ��  T     �� ���       ���� �����  �  5         ����
  G H           #uW� �     �����   p   ��  T     �� ���       ���� $�����  �  5         ����
  I J           )|_� �     ����ĸ  @�   ��  T     �� ���       ���� +�����  �  5         ����
  K L           /�g� �     ������  `�   ��  T     �� ���       ���� 3�����  �  5         ����
  M N           5�o�     ����H�  ��   ��  T	     �� ���       ���� <�����  �  5         ����
  5 6           �� �� �     ����"�  ��   ��  b      �� ���        ���� �����  �  6         ����
  7 8           �� �� �     ����Ƙ  ��   ��  b     �� ���        ���� �����  �  6         ����
  9 :           �� �� �     ����j�  6	   ��  b     �� ���        ���� �����  �  6         ����
  ; <           �� �� �     �����  �$	   ��  b     �� ���       ���� �����  �  6         ����
  = >           �� �� �     ������  n=	   ��  b     �� ���       ���� �����  �  6         ����
  ? @           �� �� �     ����V�  
V	   ��  b     �� ���       ���� �����  �  6         ����
  B C           �� �� �     ������  �n	   ��  b     �� ���       ���� �����  �  6         ����
  D E           �� �� �     ������  B�	   ��  b     �� ���       ���� �����  �  6         ����
  F G           �� �� �     ����B�  ޟ	   ��  b     �� ���       ���� &�����  �  6         ����
  H I           �� �� �     �����  z�	   ��  b	     �� ���       ���� /�����  �  6         ����
  9 :           �� �� �     ����v�  `�
   ��  c      �� ���        ���� �����  �  7         ����
  ; <           �� �� �     ����8�  ��
   ��  c     �� ���        ���� �����  �  7         ����
  = >           �� �� �     ������  ��
   ��  c     �� ���        ���� �����  �  7         ����
  ? @           �� �� �     ������  �   ��  c     �� ���       ���� �����  �  7         ����
  A B           �� �� �     ����~�  �7   ��  c     �� ���       ���� �����  �  7         ����
  C D           �� �� �     ����@�   T   ��  c     �� ���       ���� �����  �  7         ����
  F G           �� �� �     �����   p   ��  c     �� ���       ���� $�����  �  7         ����
  H I           � � �     ����ĸ  @�   ��  c     �� ���       ���� +�����  �  7         ����
  J K           � � �     ������  `�   ��  c     �� ���       ���� 3�����  �  7         ����
  L M           � � �     ����H�  ��   ��  c	     �� ���       ���� <�����  �  7         ����
  ) *           � !�� �     ����"�  ��   ��  q      �� ���        ���� �����  �  8         ����
  + ,           � '�� �     ����Ƙ  ��   ��  q     �� ���        ���� �����  �  8         ����
  - .           � -� �     ����j�  6	   ��  q     �� ���        ���� �����  �  8         ����
  / 0           � 3� �     �����  �$	   ��  q     �� ���       ���� �����  �  8         ����
  1 2           � 9� �     ������  n=	   ��  q     �� ���       ���� �����  �  8         ����
  3 4           � ?� �     ����V�  
V	   ��  q     �� ���       ���� �����  �  8         ����
  5 6           � E$� �     ������  �n	   ��  q     �� ���       ���� �����  �  8         ����
  7 8            K,� �     ������  B�	   ��  q     �� ���       ���� �����  �  8         ����
  9 :           Q4� �     ����B�  ޟ	   ��  q     �� ���       ���� &�����  �  8         ����
  ; <           W<� �     �����  z�	   ��  q	     �� ���       ���� /�����  �  8         ����
  , -           � >"� �     ����v�  `�
   ��  r      �� ���        ���� �����  �  9         ����
  . /           � E*� �     ����8�  ��
   ��  r     �� ���        ���� �����  �  9         ����
  0 1           L2� �     ������  ��
   ��  r     �� ���        ���� �����  �  9         ����
  2 3           S:� �     ������  �   ��  r     �� ���       ���� �����  �  9         ����
  4 5           ZB� �     ����~�  �7   ��  r     �� ���       ���� �����  �  9         ����
  6 7           aJ� �     ����@�   T   ��  r     �� ���       ���� �����  �  9         ����
  8 9           hR� �     �����   p   ��  r     �� ���       ���� $�����  �  9         ����
  : ;            oZ� �     ����ĸ  @�   ��  r     �� ���       ���� +�����  �  9         ����
  < =           &vb�     ������  `�   ��  r     �� ���       ���� 3�����  �  9         ����
  > ?           ,}j	�     ����H�  ��   ��  r	     �� ���       ���� <�����  �  9         ����
  8 9           ��� � �     ����"�  ��   ��  �      ��  ���        ���� �����  �  :         ����
  : ;           ��� � �     ����Ƙ  ��   ��  �     ��  ���        ���� �����  �  :         ����
  < =           ��� � �     ����j�  6	   ��  �     ��  ���        ���� �����  �  :         ����
  > ?           ��� � �     �����  �$	   ��  �     ��  ���       ���� �����  �  :         ����
  @ A           ��� � �     ������  n=	   ��  �     ��  ���       ���� �����  �  :         ����
  B C           ��� � �     ����V�  
V	   ��  �     ��  ���       ���� �����  �  :         ����
  E F           ��� � �     ������  �n	   ��  �     ��  ���       ���� �����  �  :         ����
  G H           ��� � �     ������  B�	   ��  �     ��  ���       ���� �����  �  :         ����
  I J           ��� � �     ����B�  ޟ	   ��  �     ��  ���       ���� &�����  �  :         ����
  K L           ��� � �     �����  z�	   ��  �	     ��  ���       ���� /�����  �  :         ����
  < =           ��� � �     ����v�  `�
   ��  �      ��  ���        ���� �����  �  ;         ����
  > ?           ��� � �     ����8�  ��
   ��  �     ��  ���        ���� �����  �  ;         ����
  @ A           ��� � �     ������  ��
   ��  �     ��  ���        ���� �����  �  ;         ����
  B C           ��� � �     ������  �   ��  �     ��  ���       ���� �����  �  ;         ����
  D E           ��� � �     ����~�  �7   ��  �     ��  ���       ���� �����  �  ;         ����
  F G           ��� � �     ����@�   T   ��  �     ��  ���       ���� �����  �  ;         ����
  I J           ��� � �     �����   p   ��  �     ��  ���       ���� $�����  �  ;         ����
  K L           ��� � �     ����ĸ  @�   ��  �     ��  ���       ���� +�����  �  ;         ����
  M N           ��� �     ������  `�   ��  �     ��  ���       ���� 3�����  �  ;         ����
  O P           ��� �     ����H�  ��   ��  �	     ��  ���       ���� <�����  �  ;         ����
   5 6           � !�� �     ����"�  ��   ��  �      ��! ���        ���� �����  �  <         ����
   7 8           � '�� �     ����Ƙ  ��   ��  �     ��! ���        ���� �����  �  <         ����
   9 :           � -� �     ����j�  6	   ��  �     ��! ���        ���� �����  �  <         ����
   ; <           � 3� �     �����  �$	   ��  �     ��! ���       ���� �����  �  <         ����
   = >           � 9� �     ������  n=	   ��  �     ��! ���       ���� �����  �  <         ����
   ? @           � ?� �     ����V�  
V	   ��  �     ��! ���       ���� �����  �  <         ����
   B C           � E&� �     ������  �n	   ��  �     ��! ���       ���� �����  �  <         ����
   D E           � K.� �     ������  B�	   ��  �     ��! ���       ���� �����  �  <         ����
   F G            Q6� �     ����B�  ޟ	   ��  �     ��! ���       ���� &�����  �  <         ����
   H I           W>� �     �����  z�	   ��  �	     ��! ���       ���� /�����  �  <         ����
   9 :           � >$� �     ����v�  `�
   ��  �      ��! ���        ���� �����  �  =         ����
   ; <           � E,� �     ����8�  ��
   ��  �     ��! ���        ���� �����  �  =         ����
   = >           � L4� �     ������  ��
   ��  �     ��! ���        ���� �����  �  =         ����
   ? @           S<� �     ������  �   ��  �     ��! ���       ���� �����  �  =         ����
   A B           ZD� �     ����~�  �7   ��  �     ��! ���       ���� �����  �  =         ����
   C D           aL� �     ����@�   T   ��  �     ��! ���       ���� �����  �  =         ����
   F G           hT� �     �����   p   ��  �     ��! ���       ���� $�����  �  =         ����
   H I           o\� �     ����ĸ  @�   ��  �     ��! ���       ���� +�����  �  =         ����
   J K            vd� �     ������  `�   ��  �     ��! ���       ���� 3�����  �  =         ����
   L M           &}l� �     ����H�  ��   ��  �	     ��! ���       ���� <�����  �  =         ����  F G           5� � �     ������  �<   ��  �      �� ���        ���� �����  �  >         ����  H I           <� � �     ����:�  fU   ��  �     �� ���        ���� �����  �  >         ����  J K           C� � �     ����ޏ  n   ��  �     �� ���        ���� �����  �  >         ����  M N           %J� � �     ������  ��   ��  �     �� ���       ���� �����  �  >         ����  O P           -Q� � �     ����&�  :�   ��  �     �� ���       ���� �����  �  >         ����  Q R           5X� � �     ����ʔ  ַ   ��  �     �� ���       ���� �����  �  >         ����  S T           =_� � �     ����n�  r�   ��  �     �� ���       ���� �����  �  >         ����  U V           Ef� � �     �����  �   ��  �     �� ���       ���� �����  �  >         ����  X Y           Mm� � �     ������  �	   ��  �     �� ���       ���� &�����  �  >         ����  Z [           Ut� � �     ����Z�  F	   ��  �	     �� ���       ���� /�����  �  >         ����  K L           ;[� � �     �����  �
   ��  �      �� ���        ���� �����  �  ?         ����  M N           Cb� � �     ������  �:
   ��  �     �� ���        ���� �����  �  ?         ����  O P           Ki� � �     ����n�  �V
   ��  �     �� ���        ���� �����  �  ?         ����  R S           Sp� � �     ����0�   s
   ��  �     �� ���       ���� �����  �  ?         ����  T U           [w� � �     �����   �
   ��  �     �� ���       ���� �����  �  ?         ����  V W           c~� � �     ������  @�
   ��  �     �� ���       ���� �����  �  ?         ����  X Y           k�� � �     ����v�  `�
   ��  �     �� ���       ���� $�����  �  ?         ����  Z [           s�� � �     ����8�  ��
   ��  �     �� ���       ���� +�����  �  ?         ����  ] ^           {�� �     ������  ��
   ��  �     �� ���       ���� 3�����  �  ?         ����  _ `           ��� �     ������  �   ��  �	     �� ���       ���� <�����  �  ?         ����  7 8           � ;� �     ������  �<   ��  �      �� ���        ���� �����  �  @         ����  9 :           � A� �     ����:�  fU   ��  �     �� ���        ���� �����  �  @         ����  ; <           � G� �     ����ޏ  n   ��  �     �� ���        ���� �����  �  @         ����  = >           � M� �     ������  ��   ��  �     �� ���       ���� �����  �  @         ����  ? @           S&� �     ����&�  :�   ��  �     �� ���       ���� �����  �  @         ����  A B           	Y.� �     ����ʔ  ַ   ��  �     �� ���       ���� �����  �  @         ����  D E           _6� �     ����n�  r�   ��  �     �� ���       ���� �����  �  @         ����  F G           e>� �     �����  �   ��  �     �� ���       ���� �����  �  @         ����  H I           kF� �     ������  �	   ��  �     �� ���       ���� &�����  �  @         ����  J K           !qN� �     ����Z�  F	   ��  �	     �� ���       ���� /�����  �  @         ����  ; <           X4� �     �����  �
   ��  �      �� ���        ���� �����  �  A         ����  = >           _<� �     ������  �:
   ��  �     �� ���        ���� �����  �  A         ����  ? @           fD� �     ����n�  �V
   ��  �     �� ���        ���� �����  �  A         ����  A B           mL� �     ����0�   s
   ��  �     �� ���       ���� �����  �  A         ����  C D           #tT� �     �����   �
   ��  �     �� ���       ���� �����  �  A         ����  E F           ){\� �     ������  @�
   ��  �     �� ���       ���� �����  �  A         ����  H I           /�d� �     ����v�  `�
   ��  �     �� ���       ���� $�����  �  A         ����  J K           5�l� �     ����8�  ��
   ��  �     �� ���       ���� +�����  �  A         ����  L M           ;�t� �     ������  ��
   ��  �     �� ���       ���� 3�����  �  A         ����  N O           A�|�     ������  �   ��  �	     �� ���       ���� <�����  �  A         ����  6 7           �� �� �     ������  �<   ��  �      �� ���        ���� �����  �  B         ����  8 9           �� �� �     ����:�  fU   ��  �     �� ���        ���� �����  �  B         ����  : ;           �� �� �     ����ޏ  n   ��  �     �� ���        ���� �����  �  B         ����  < =           �� �� �     ������  ��   ��  �     �� ���       ���� �����  �  B         ����  > ?           �� �� �     ����&�  :�   ��  �     �� ���       ���� �����  �  B         ����  @ A           �� �� �     ����ʔ  ַ   ��  �     �� ���       ���� �����  �  B         ����  C D           �� �� �     ����n�  r�   ��  �     �� ���       ���� �����  �  B         ����  E F           �� �� �     �����  �   ��  �     �� ���       ���� �����  �  B         ����  G H           �� �� �     ������  �	   ��  �     �� ���       ���� &�����  �  B         ����  I J           �� �� �     ����Z�  F	   ��  �	     �� ���       ���� /�����  �  B         ����  : ;           �� �� �     �����  �
   ��  �      �� ���        ���� �����  �  C         ����  < =           �� �� �     ������  �:
   ��  �     �� ���        ���� �����  �  C         ����  > ?           �� �� �     ����n�  �V
   ��  �     �� ���        ���� �����  �  C         ����  @ A           �� �� �     ����0�   s
   ��  �     �� ���       ���� �����  �  C         ����  B C           �� �� �     �����   �
   ��  �     �� ���       ���� �����  �  C         ����  D E           � � �     ������  @�
   ��  �     �� ���       ���� �����  �  C         ����  G H           	� 	� �     ����v�  `�
   ��  �     �� ���       ���� $�����  �  C         ����  I J           � � �     ����8�  ��
   ��  �     �� ���       ���� +�����  �  C         ����  K L           � � �     ������  ��
   ��  �     �� ���       ���� 3�����  �  C         ����  M N           !� !� �     ������  �   ��  �	     �� ���       ���� <�����  �  C         ����  ) *           � *�� �     ������  �<   ��  �      �� ���        ���� �����  �  D         ����  + ,           � 0� �     ����:�  fU   ��  �     �� ���        ���� �����  �  D         ����  - .           � 6� �     ����ޏ  n   ��  �     �� ���        ���� �����  �  D         ����  / 0           � <� �     ������  ��   ��  �     �� ���       ���� �����  �  D         ����  1 2           � B� �     ����&�  :�   ��  �     �� ���       ���� �����  �  D         ����  3 4           � H%� �     ����ʔ  ַ   ��  �     �� ���       ���� �����  �  D         ����  5 6            N-� �     ����n�  r�   ��  �     �� ���       ���� �����  �  D         ����  7 8           T5� �     �����  �   ��  �     �� ���       ���� �����  �  D         ����  9 :           Z=� �     ������  �	   ��  �     �� ���       ���� &�����  �  D         ����  ; <           `E� �     ����Z�  F	   ��  �	     �� ���       ���� /�����  �  D         ����  , -           � G+� �     �����  �
   ��  �      �� ���        ���� �����  �  E         ����  . /           N3� �     ������  �:
   ��  �     �� ���        ���� �����  �  E         ����  0 1           U;� �     ����n�  �V
   ��  �     �� ���        ���� �����  �  E         ����  2 3           \C� �     ����0�   s
   ��  �     �� ���       ���� �����  �  E         ����  4 5           cK� �     �����   �
   ��  �     �� ���       ���� �����  �  E         ����  6 7           jS �     ������  @�
   ��  �     �� ���       ���� �����  �  E         ����  8 9            q[�     ����v�  `�
   ��  �     �� ���       ���� $�����  �  E         ����  : ;           &xc�     ����8�  ��
   ��  �     �� ���       ���� +�����  �  E         ����  < =           ,k�     ������  ��
   ��  �     �� ���       ���� 3�����  �  E         ����  > ?           2�s�     ������  �   ��  �	     �� ���       ���� <�����  �  E         ����  9 :           ��� � �     ������  �<   ��  �      ��  ���        ���� �����  �  F         ����  ; <           ��� � �     ����:�  fU   ��  �     ��  ���        ���� �����  �  F         ����  = >           ��� � �     ����ޏ  n   ��  �     ��  ���        ���� �����  �  F         ����  ? @           ��� � �     ������  ��   ��  �     ��  ���       ���� �����  �  F         ����  A B           ��� � �     ����&�  :�   ��  �     ��  ���       ���� �����  �  F         ����  C D           ��� � �     ����ʔ  ַ   ��  �     ��  ���       ���� �����  �  F         ����  F G           ��� � �     ����n�  r�   ��  �     ��  ���       ���� �����  �  F         ����  H I           ��� � �     �����  �   ��  �     ��  ���       ���� �����  �  F         ����  J K           ��� � �     ������  �	   ��  �     ��  ���       ���� &�����  �  F         ����  L M           ��� � �     ����Z�  F	   ��  �	     ��  ���       ���� /�����  �  F         ����  = >           ��� � �     �����  �
   ��  �      ��  ���        ���� �����  �  G         ����  ? @           ��� � �     ������  �:
   ��  �     ��  ���        ���� �����  �  G         ����  A B           ��� � �     ����n�  �V
   ��  �     ��  ���        ���� �����  �  G         ����  C D           ��� � �     ����0�   s
   ��  �     ��  ���       ���� �����  �  G         ����  E F           ��� � �     �����   �
   ��  �     ��  ���       ���� �����  �  G         ����  G H           ��� � �     ������  @�
   ��  �     ��  ���       ���� �����  �  G         ����  J K           ��� � �     ����v�  `�
   ��  �     ��  ���       ���� $�����  �  G         ����  L M           ��� � �     ����8�  ��
   ��  �     ��  ���       ���� +�����  �  G         ����  N O           ��� �     ������  ��
   ��  �     ��  ���       ���� 3�����  �  G         ����  P Q           �� �     ������  �   ��  �	     ��  ���       ���� <�����  �  G         ����   6 7           � !�� �     ������  �<   ��  �      ��! ���        ���� �����  �  H         ����   8 9           � '� �     ����:�  fU   ��  �     ��! ���        ���� �����  �  H         ����   : ;           � -� �     ����ޏ  n   ��  �     ��! ���        ���� �����  �  H         ����   < =           � 3� �     ������  ��   ��  �     ��! ���       ���� �����  �  H         ����   > ?           � 9� �     ����&�  :�   ��  �     ��! ���       ���� �����  �  H         ����   @ A           � ?&� �     ����ʔ  ַ   ��  �     ��! ���       ���� �����  �  H         ����   C D           � E.� �     ����n�  r�   ��  �     ��! ���       ���� �����  �  H         ����   E F           � K6� �     �����  �   ��  �     ��! ���       ���� �����  �  H         ����   G H            Q>� �     ������  �	   ��  �     ��! ���       ���� &�����  �  H         ����   I J           WF� �     ����Z�  F	   ��  �	     ��! ���       ���� /�����  �  H         ����   : ;           � >,� �     �����  �
   ��  �      ��! ���        ���� �����  �  I         ����   < =           � E4� �     ������  �:
   ��  �     ��! ���        ���� �����  �  I         ����   > ?           � L<� �     ����n�  �V
   ��  �     ��! ���        ���� �����  �  I         ����   @ A           SD� �     ����0�   s
   ��  �     ��! ���       ���� �����  �  I         ����   B C           ZL� �     �����   �
   ��  �     ��! ���       ���� �����  �  I         ����   D E           aT� �     ������  @�
   ��  �     ��! ���       ���� �����  �  I         ����   G H           h\� �     ����v�  `�
   ��  �     ��! ���       ���� $�����  �  I         ����   I J           od� �     ����8�  ��
   ��  �     ��! ���       ���� +�����  �  I         ����   K L            vl� �     ������  ��
   ��  �     ��! ���       ���� 3�����  �  I         ����   M N           &}t� �     ������  �   ��  �	     ��! ���       ���� <�����  �  I         ����  G H           5� � �     ����B�  �		   ��  �      �� ���        ���� �����  �  J         ����  I J           "<� � �     �����  z"	   ��  �     �� ���        ���� �����  �  J         ����  K L           *C� � �     ������  ;	   ��  �     �� ���        ���� �����  �  J         ����  N O           2J� � �     ����.�  �S	   ��  �     �� ���       ���� �����  �  J         ����  P Q           :Q� � �     ����Ҡ  Nl	   ��  �     �� ���       ���� �����  �  J         ����  R S           BX� � �     ����v�  �	   ��  �     �� ���       ���� �����  �  J         ����  T U           J_� � �     �����  ��	   ��  �     �� ���       ���� �����  �  J         ����  V W           Rf� � �     ������  "�	   ��  �     �� ���       ���� �����  �  J         ����  Y Z           Zm� � �     ����b�  ��	   ��  �     �� ���       ���� &�����  �  J         ����  [ \           bt� � �     �����  Z�	   ��  �	     �� ���       ���� /�����  �  J         ����  L M           H[� � �     ������  `�
   ��  �      �� ���        ���� �����  �  K         ����  N O           Pb� � �     ����X�  �   ��  �     �� ���        ���� �����  �  K         ����  P Q           Xi� � �     �����  �1   ��  �     �� ���        ���� �����  �  K         ����  S T           `p� � �     ����ܴ  �M   ��  �     �� ���       ���� �����  �  K         ����  U V           hw� � �     ������  �i   ��  �     �� ���       ���� �����  �  K         ����  W X           p~� � �     ����`�   �   ��  �     �� ���       ���� �����  �  K         ����  Y Z           x�� � �     ����"�   �   ��  �     �� ���       ���� $�����  �  K         ����  [ \           ��� � �     �����  @�   ��  �     �� ���       ���� +�����  �  K         ����  ^ _           ��� �     ������  `�   ��  �     �� ���       ���� 3�����  �  K         ����  ` a           ��� �     ����h�  ��   ��  �	     �� ���       ���� <�����  �  K         ����  7 8           � H� �     ����B�  �		   ��        �� ���        ���� �����  �  L         ����  9 :           � N� �     �����  z"	   ��       �� ���        ���� �����  �  L         ����  ; <           T#� �     ������  ;	   ��       �� ���        ���� �����  �  L         ����  = >           
Z+� �     ����.�  �S	   ��       �� ���       ���� �����  �  L         ����  ? @           `3� �     ����Ҡ  Nl	   ��       �� ���       ���� �����  �  L         ����  A B           f;� �     ����v�  �	   ��       �� ���       ���� �����  �  L         ����  D E           lC� �     �����  ��	   ��       �� ���       ���� �����  �  L         ����  F G           "rK� �     ������  "�	   ��       �� ���       ���� �����  �  L         ����  H I           (xS� �     ����b�  ��	   ��       �� ���       ���� &�����  �  L         ����  J K           .~[� �     �����  Z�	   ��  	     �� ���       ���� /�����  �  L         ����  ; <           eA� �     ������  `�
   ��        �� ���        ���� �����  �  M         ����  = >           lI� �     ����X�  �   ��       �� ���        ���� �����  �  M         ����  ? @           $sQ� �     �����  �1   ��       �� ���        ���� �����  �  M         ����  A B           *zY� �     ����ܴ  �M   ��       �� ���       ���� �����  �  M         ����  C D           0�a� �     ������  �i   ��       �� ���       ���� �����  �  M         ����  E F           6�i� �     ����`�   �   ��       �� ���       ���� �����  �  M         ����  H I           <�q� �     ����"�   �   ��       �� ���       ���� $�����  �  M         ����  J K           B�y� �     �����  @�   ��       �� ���       ���� +�����  �  M         ����  L M           H��� �     ������  `�   ��       �� ���       ���� 3�����  �  M         ����  N O           N���     ����h�  ��   ��  	     �� ���       ���� <�����  �  M         ����  6 7           �� �� �     ����B�  �		   ��        �� ���        ���� �����  �  N         ����  8 9           �� �� �     �����  z"	   ��       �� ���        ���� �����  �  N         ����  : ;           �� �� �     ������  ;	   ��       �� ���        ���� �����  �  N         ����  < =           �� �� �     ����.�  �S	   ��       �� ���       ���� �����  �  N         ����  > ?           �� �� �     ����Ҡ  Nl	   ��       �� ���       ���� �����  �  N         ����  @ A           �� �� �     ����v�  �	   ��       �� ���       ���� �����  �  N         ����  C D           �� �� �     �����  ��	   ��       �� ���       ���� �����  �  N         ����  E F           �� �� �     ������  "�	   ��       �� ���       ���� �����  �  N         ����  G H           �� �� �     ����b�  ��	   ��       �� ���       ���� &�����  �  N         ����  I J           �� �� �     �����  Z�	   ��  	     �� ���       ���� /�����  �  N         ����  : ;           �� �� �     ������  `�
   ��        �� ���        ���� �����  �  O         ����  < =           �� �� �     ����X�  �   ��       �� ���        ���� �����  �  O         ����  > ?           �� �� �     �����  �1   ��       �� ���        ���� �����  �  O         ����  @ A           �� �� �     ����ܴ  �M   ��       �� ���       ���� �����  �  O         ����  B C           � � �     ������  �i   ��       �� ���       ���� �����  �  O         ����  D E           � � �     ����`�   �   ��       �� ���       ���� �����  �  O         ����  G H           � � �     ����"�   �   ��       �� ���       ���� $�����  �  O         ����  I J           � � �     �����  @�   ��       �� ���       ���� +�����  �  O         ����  K L           &� &� �     ������  `�   ��       �� ���       ���� 3�����  �  O         ����  M N           .� .� �     ����h�  ��   ��  	     �� ���       ���� <�����  �  O         ����  ) *           � 3� �     ����B�  �		   ��  %      �� ���        ���� �����  �  P         ����  + ,           � 9� �     �����  z"	   ��  %     �� ���        ���� �����  �  P         ����  - .           � ?� �     ������  ;	   ��  %     �� ���        ���� �����  �  P         ����  / 0           � E� �     ����.�  �S	   ��  %     �� ���       ���� �����  �  P         ����  1 2           � K&� �     ����Ҡ  Nl	   ��  %     �� ���       ���� �����  �  P         ����  3 4           � Q.� �     ����v�  �	   ��  %     �� ���       ���� �����  �  P         ����  5 6           W6� �     �����  ��	   ��  %     �� ���       ���� �����  �  P         ����  7 8           ]>� �     ������  "�	   ��  %     �� ���       ���� �����  �  P         ����  9 :           cF� �     ����b�  ��	   ��  %     �� ���       ���� &�����  �  P         ����  ; <           iN� �     �����  Z�	   ��  %	     �� ���       ���� /�����  �  P         ����  , -           P4� �     ������  `�
   ��  &      �� ���        ���� �����  �  Q         ����  . /           W<� �     ����X�  �   ��  &     �� ���        ���� �����  �  Q         ����  0 1           ^D� �     �����  �1   ��  &     �� ���        ���� �����  �  Q         ����  2 3           eL� �     ����ܴ  �M   ��  &     �� ���       ���� �����  �  Q         ����  4 5           lT� �     ������  �i   ��  &     �� ���       ���� �����  �  Q         ����  6 7           s\�     ����`�   �   ��  &     �� ���       ���� �����  �  Q         ����  8 9           %zd�     ����"�   �   ��  &     �� ���       ���� $�����  �  Q         ����  : ;           +�l�     �����  @�   ��  &     �� ���       ���� +�����  �  Q         ����  < =           1�t�     ������  `�   ��  &     �� ���       ���� 3�����  �  Q         ����  > ?           7�|�     ����h�  ��   ��  &	     �� ���       ���� <�����  �  Q         ����  9 :           ��� � �     ����B�  �		   ��  4      ��  ���        ���� �����  �  R         ����  ; <           ��� � �     �����  z"	   ��  4     ��  ���        ���� �����  �  R         ����  = >           ��� � �     ������  ;	   ��  4     ��  ���        ���� �����  �  R         ����  ? @           ��� � �     ����.�  �S	   ��  4     ��  ���       ���� �����  �  R         ����  A B           ��� � �     ����Ҡ  Nl	   ��  4     ��  ���       ���� �����  �  R         ����  C D           ��� � �     ����v�  �	   ��  4     ��  ���       ���� �����  �  R         ����  F G           ��� � �     �����  ��	   ��  4     ��  ���       ���� �����  �  R         ����  H I           ��� � �     ������  "�	   ��  4     ��  ���       ���� �����  �  R         ����  J K           ��� � �     ����b�  ��	   ��  4     ��  ���       ���� &�����  �  R         ����  L M           ��� � �     �����  Z�	   ��  4	     ��  ���       ���� /�����  �  R         ����  = >           ��� � �     ������  `�
   ��  5      ��  ���        ���� �����  �  S         ����  ? @           ��� � �     ����X�  �   ��  5     ��  ���        ���� �����  �  S         ����  A B           ��� � �     �����  �1   ��  5     ��  ���        ���� �����  �  S         ����  C D           ��� � �     ����ܴ  �M   ��  5     ��  ���       ���� �����  �  S         ����  E F           ��� � �     ������  �i   ��  5     ��  ���       ���� �����  �  S         ����  G H           ��� � �     ����`�   �   ��  5     ��  ���       ���� �����  �  S         ����  J K           ��� � �     ����"�   �   ��  5     ��  ���       ���� $�����  �  S         ����  L M           ��� � �     �����  @�   ��  5     ��  ���       ���� +�����  �  S         ����  N O           �� �     ������  `�   ��  5     ��  ���       ���� 3�����  �  S         ����  P Q           �� �     ����h�  ��   ��  5	     ��  ���       ���� <�����  �  S         ����   6 7           � !� �     ����B�  �		   ��  C      ��! ���        ���� �����  �  T         ����   8 9           � '� �     �����  z"	   ��  C     ��! ���        ���� �����  �  T         ����   : ;           � -� �     ������  ;	   ��  C     ��! ���        ���� �����  �  T         ����   < =           � 3� �     ����.�  �S	   ��  C     ��! ���       ���� �����  �  T         ����   > ?           � 9&� �     ����Ҡ  Nl	   ��  C     ��! ���       ���� �����  �  T         ����   @ A           � ?.� �     ����v�  �	   ��  C     ��! ���       ���� �����  �  T         ����   C D           � E6� �     �����  ��	   ��  C     ��! ���       ���� �����  �  T         ����   E F           � K>� �     ������  "�	   ��  C     ��! ���       ���� �����  �  T         ����   G H            QF� �     ����b�  ��	   ��  C     ��! ���       ���� &�����  �  T         ����   I J           WN� �     �����  Z�	   ��  C	     ��! ���       ���� /�����  �  T         ����   : ;           � >4� �     ������  `�
   ��  D      ��! ���        ���� �����  �  U         ����   < =           � E<� �     ����X�  �   ��  D     ��! ���        ���� �����  �  U         ����   > ?           � LD� �     �����  �1   ��  D     ��! ���        ���� �����  �  U         ����   @ A           SL� �     ����ܴ  �M   ��  D     ��! ���       ���� �����  �  U         ����   B C           ZT� �     ������  �i   ��  D     ��! ���       ���� �����  �  U         ����   D E           a\� �     ����`�   �   ��  D     ��! ���       ���� �����  �  U         ����   G H           hd� �     ����"�   �   ��  D     ��! ���       ���� $�����  �  U         ����   I J           ol� �     �����  @�   ��  D     ��! ���       ���� +�����  �  U         ����   K L            vt� �     ������  `�   ��  D     ��! ���       ���� 3�����  �  U         ����   M N           &}|� �     ����h�  ��   ��  D	     ��! ���       ���� <�����  �  U         ����  G H           5� � �     ����қ  N!	   ��  R      �� ���        ���� �����  �  V         ����  I J           %<� � �     ����v�  �9	   ��  R     �� ���        ���� �����  �  V         ����  K L           -C� � �     �����  �R	   ��  R     �� ���        ���� �����  �  V         ����  N O           5J� � �     ������  "k	   ��  R     �� ���       ���� �����  �  V         ����  P Q           =Q� � �     ����b�  ��	   ��  R     �� ���       ���� �����  �  V         ����  R S           EX� � �     �����  Z�	   ��  R     �� ���       ���� �����  �  V         ����  T U           M_� � �     ������  ��	   ��  R     �� ���       ���� �����  �  V         ����  V W           Uf� � �     ����N�  ��	   ��  R     �� ���       ���� �����  �  V         ����  Y Z           ]m� � �     �����  .�	   ��  R     �� ���       ���� &�����  �  V         ����  [ \           et� � �     ������  ��	   ��  R	     �� ���       ���� /�����  �  V         ����  L M           K[� � �     ����&�  `   ��  S      �� ���        ���� �����  �  W         ����  N O           Sb� � �     �����  �.   ��  S     �� ���        ���� �����  �  W         ����  P Q           [i� � �     ������  �J   ��  S     �� ���        ���� �����  �  W         ����  S T           cp� � �     ����l�  �f   ��  S     �� ���       ���� �����  �  W         ����  U V           kw� � �     ����.�  ��   ��  S     �� ���       ���� �����  �  W         ����  W X           s~� � �     �����   �   ��  S     �� ���       ���� �����  �  W         ����  Y Z           {�� � �     ������   �   ��  S     �� ���       ���� $�����  �  W         ����  [ \           ��� � �     ����t�  @�   ��  S     �� ���       ���� +�����  �  W         ����  ^ _           ��� �     ����6�  `�   ��  S     �� ���       ���� 3�����  �  W         ����  ` a           ��� �     ������  �   ��  S	     �� ���       ���� <�����  �  W         ����  7 8           � K� �     ����қ  N!	   ��  a      �� ���        ���� �����  �  X         ����  9 :           Q� �     ����v�  �9	   ��  a     �� ���        ���� �����  �  X         ����  ; <           W&� �     �����  �R	   ��  a     �� ���        ���� �����  �  X         ����  = >           ].� �     ������  "k	   ��  a     �� ���       ���� �����  �  X         ����  ? @           c6� �     ����b�  ��	   ��  a     �� ���       ���� �����  �  X         ����  A B           i>� �     �����  Z�	   ��  a     �� ���       ���� �����  �  X         ����  D E           oF� �     ������  ��	   ��  a     �� ���       ���� �����  �  X         ����  F G           %uN� �     ����N�  ��	   ��  a     �� ���       ���� �����  �  X         ����  H I           +{V� �     �����  .�	   ��  a     �� ���       ���� &�����  �  X         ����  J K           1�^� �     ������  ��	   ��  a	     �� ���       ���� /�����  �  X         ����  ; <           hD� �     ����&�  `   ��  b      �� ���        ���� �����  �  Y         ����  = >           !oL� �     �����  �.   ��  b     �� ���        ���� �����  �  Y         ����  ? @           'vT� �     ������  �J   ��  b     �� ���        ���� �����  �  Y         ����  A B           -}\� �     ����l�  �f   ��  b     �� ���       ���� �����  �  Y         ����  C D           3�d� �     ����.�  ��   ��  b     �� ���       ���� �����  �  Y         ����  E F           9�l� �     �����   �   ��  b     �� ���       ���� �����  �  Y         ����  H I           ?�t� �     ������   �   ��  b     �� ���       ���� $�����  �  Y         ����  J K           E�|� �     ����t�  @�   ��  b     �� ���       ���� +�����  �  Y         ����  L M           K��� �     ����6�  `�   ��  b     �� ���       ���� 3�����  �  Y         ����  N O           Q���     ������  �   ��  b	     �� ���       ���� <�����  �  Y         ����  6 7           �� �� �     ����қ  N!	   ��  p      �� ���        ���� �����  �  Z         ����  8 9           �� �� �     ����v�  �9	   ��  p     �� ���        ���� �����  �  Z         ����  : ;           �� �� �     �����  �R	   ��  p     �� ���        ���� �����  �  Z         ����  < =           �� �� �     ������  "k	   ��  p     �� ���       ���� �����  �  Z         ����  > ?           �� �� �     ����b�  ��	   ��  p     �� ���       ���� �����  �  Z         ����  @ A           �� �� �     �����  Z�	   ��  p     �� ���       ���� �����  �  Z         ����  C D           �� �� �     ������  ��	   ��  p     �� ���       ���� �����  �  Z         ����  E F           �� �� �     ����N�  ��	   ��  p     �� ���       ���� �����  �  Z         ����  G H           �� �� �     �����  .�	   ��  p     �� ���       ���� &�����  �  Z         ����  I J           � � �     ������  ��	   ��  p	     �� ���       ���� /�����  �  Z         ����  : ;           �� �� �     ����&�  `   ��  q      �� ���        ���� �����  �  [         ����  < =           �� �� �     �����  �.   ��  q     �� ���        ���� �����  �  [         ����  > ?           �� �� �     ������  �J   ��  q     �� ���        ���� �����  �  [         ����  @ A           � � �     ����l�  �f   ��  q     �� ���       ���� �����  �  [         ����  B C           	� 	� �     ����.�  ��   ��  q     �� ���       ���� �����  �  [         ����  D E           � � �     �����   �   ��  q     �� ���       ���� �����  �  [         ����  G H           � � �     ������   �   ��  q     �� ���       ���� $�����  �  [         ����  I J           !� !� �     ����t�  @�   ��  q     �� ���       ���� +�����  �  [         ����  K L           )� )� �     ����6�  `�   ��  q     �� ���       ���� 3�����  �  [         ����  M N           1� 1� �     ������  �   ��  q	     �� ���       ���� <�����  �  [         ����  ) *           � 6	� �     ����қ  N!	   ��        �� ���        ���� �����  �  \         ����  + ,           � <� �     ����v�  �9	   ��       �� ���        ���� �����  �  \         ����  - .           � B� �     �����  �R	   ��       �� ���        ���� �����  �  \         ����  / 0           � H!� �     ������  "k	   ��       �� ���       ���� �����  �  \         ����  1 2           N)� �     ����b�  ��	   ��       �� ���       ���� �����  �  \         ����  3 4           	T1� �     �����  Z�	   ��       �� ���       ���� �����  �  \         ����  5 6           Z9� �     ������  ��	   ��       �� ���       ���� �����  �  \         ����  7 8           `A� �     ����N�  ��	   ��       �� ���       ���� �����  �  \         ����  9 :           fI� �     �����  .�	   ��       �� ���       ���� &�����  �  \         ����  ; <           !lQ� �     ������  ��	   ��  	     �� ���       ���� /�����  �  \         ����  , -           S7� �     ����&�  `   ��  �      �� ���        ���� �����  �  ]         ����  . /           Z?� �     �����  �.   ��  �     �� ���        ���� �����  �  ]         ����  0 1           aG� �     ������  �J   ��  �     �� ���        ���� �����  �  ]         ����  2 3           hO� �     ����l�  �f   ��  �     �� ���       ���� �����  �  ]         ����  4 5           #oW �     ����.�  ��   ��  �     �� ���       ���� �����  �  ]         ����  6 7           )v_�     �����   �   ��  �     �� ���       ���� �����  �  ]         ����  8 9           /}g�     ������   �   ��  �     �� ���       ���� $�����  �  ]         ����  : ;           5�o�     ����t�  @�   ��  �     �� ���       ���� +�����  �  ]         ����  < =           ;�w�     ����6�  `�   ��  �     �� ���       ���� 3�����  �  ]         ����  > ?           A��     ������  �   ��  �	     �� ���       ���� <�����  �  ]         ����  9 :           ��� � �     ����қ  N!	   ��  �      ��  ���        ���� �����  �  ^         ����  ; <           ��� � �     ����v�  �9	   ��  �     ��  ���        ���� �����  �  ^         ����  = >           ��� � �     �����  �R	   ��  �     ��  ���        ���� �����  �  ^         ����  ? @           ��� � �     ������  "k	   ��  �     ��  ���       ���� �����  �  ^         ����  A B           ��� � �     ����b�  ��	   ��  �     ��  ���       ���� �����  �  ^         ����  C D           ��� � �     �����  Z�	   ��  �     ��  ���       ���� �����  �  ^         ����  F G           ��� � �     ������  ��	   ��  �     ��  ���       ���� �����  �  ^         ����  H I           ��� � �     ����N�  ��	   ��  �     ��  ���       ���� �����  �  ^         ����  J K           ��� � �     �����  .�	   ��  �     ��  ���       ���� &�����  �  ^         ����  L M           ��� � �     ������  ��	   ��  �	     ��  ���       ���� /�����  �  ^         ����  = >           ��� � �     ����&�  `   ��  �      ��  ���        ���� �����  �  _         ����  ? @           ��� � �     �����  �.   ��  �     ��  ���        ���� �����  �  _         ����  A B           ��� � �     ������  �J   ��  �     ��  ���        ���� �����  �  _         ����  C D           ��� � �     ����l�  �f   ��  �     ��  ���       ���� �����  �  _         ����  E F           ��� � �     ����.�  ��   ��  �     ��  ���       ���� �����  �  _         ����  G H           ��� � �     �����   �   ��  �     ��  ���       ���� �����  �  _         ����  J K           ��� � �     ������   �   ��  �     ��  ���       ���� $�����  �  _         ����  L M           � � � �     ����t�  @�   ��  �     ��  ���       ���� +�����  �  _         ����  N O           �� �     ����6�  `�   ��  �     ��  ���       ���� 3�����  �  _         ����  P Q           �� �     ������  �   ��  �	     ��  ���       ���� <�����  �  _         ����   6 7           � <� �     ����қ  N!	   ��  �      ��! ���        ���� �����  �  `         ����   8 9           � D� �     ����v�  �9	   ��  �     ��! ���        ���� �����  �  `         ����   : ;           � #L� �     �����  �R	   ��  �     ��! ���        ���� �����  �  `         ����   < =           � )T� �     ������  "k	   ��  �     ��! ���       ���� �����  �  `         ����   > ?           � /\� �     ����b�  ��	   ��  �     ��! ���       ���� �����  �  `         ����   @ A           � 5d� �     �����  Z�	   ��  �     ��! ���       ���� �����  �  `         ����   C D           � ;l� �     ������  ��	   ��  �     ��! ���       ���� �����  �  `         ����   E F           � At� �     ����N�  ��	   ��  �     ��! ���       ���� �����  �  `         ����   G H           � G|� �     �����  .�	   ��  �     ��! ���       ���� &�����  �  `         ����   I J           � M�� �     ������  ��	   ��  �	     ��! ���       ���� /�����  �  `         ����   : ;           � 3p� �     ����&�  `   ��  �      ��! ���        ���� �����  �  a         ����   < =           � :x� �     �����  �.   ��  �     ��! ���        ���� �����  �  a         ����   > ?           � A�� �     ������  �J   ��  �     ��! ���        ���� �����  �  a         ����   @ A           � H�� �     ����l�  �f   ��  �     ��! ���       ���� �����  �  a         ����   B C           � O�� �     ����.�  ��   ��  �     ��! ���       ���� �����  �  a         ����   D E           � V�� �     �����   �   ��  �     ��! ���       ���� �����  �  a         ����   G H           � ]�� �     ������   �   ��  �     ��! ���       ���� $�����  �  a         ����   I J           � d�� �     ����t�  @�   ��  �     ��! ���       ���� +�����  �  a         ����   K L           � k�� �     ����6�  `�   ��  �     ��! ���       ���� 3�����  �  a         ����   M N           � r�� �     ������  �   ��  �	     ��! ���       ���� <�����  �  a          ��� ��                        ����    �  �     �  d   �� ���        ������  ����������������        ��� ��                        ����    �  �     �  d   �� ���        ������  ����������������        ��� ��                        ����    �  �     �  d   �� ���        ������  ����������������        ��� ��                       ����    �  �     �  e   �� ���        ������  ����������������        ��� ��#    Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    Z  
                  ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    �  
                  ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��#    �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   Z  
                  ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   Z                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   �  
                  ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��# (   �                    ����    �  �     �  f   �� ���        ������  ����������������        ��� ��$    Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    Z  
                  ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    �  
                  ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$    �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   Z  
                  ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   Z                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   �  
                  ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��$ (   �                    ����    �  �     �  g   �� ���        ������  ����������������        ��� ��&    <                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    <  
                  ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    <                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    <                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    x                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    x  
                  ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    x                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��&    x                    ����    �  �     �  h   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    Z  
                  ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    �  
                  ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   Z  
                  ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   �  
                  ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  i   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    Z  
                  ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    �  
                  ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   Z  
                  ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   �  
                  ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  j   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    Z  
                  ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    �  
                  ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   Z  
                  ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   �  
                  ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �     �  k   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    Z  
                  ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    Z                    ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    �  
                  ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  l   �� ���        ������  ����������������        ��� ��    �                    ����    �  �     �  l   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �     �  l   �� ���        ������  ����������������        ��� �� (   Z  
                  ����    �  �     �  l   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �        l   �� ���        ������  ����������������        ��� �� (   Z                    ����    �  �       l   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �       l   �� ���        ������  ����������������        ��� �� (   �  
                  ����    �  �       l   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �       l   �� ���        ������  ����������������        ��� �� (   �                    ����    �  �       l   �� ���        ������  ����������������        ��� �� 
   <                    ����    �  �       m   �� ���        ������  ����������������        ��� �� 
   <  
                  ����    �  �       m   �� ���        ������  ����������������        ��� �� 
   <                    ����    �  �       m   �� ���        ������  ����������������        ��� �� 
   <                    ����    �  �     	  m   �� ���        ������  ����������������        ��� �� 
   x                    ����    �  �     
  m   �� ���        ������  ����������������        ��� �� 
   x  
                  ����    �  �       m   �� ���        ������  ����������������        ��� �� 
   x                    ����    �  �       m   �� ���        ������  ����������������        ��� �� 
   x                    ����    �  �       m   �� ���        ������  ����������������        ��� ��! 
   <                    ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   <  
                  ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   <                    ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   <                    ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   x                    ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   x  
                  ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   x                    ����    �  �       n   �� ���        ������  ����������������        ��� ��! 
   x                    ����    �  �       n   �� ���        ������  ����������������        ��� ��    <                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    <  
                  ����    �  �       o   �� ���        ������  ����������������        ��� ��    <                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    <                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    x                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    x  
                  ����    �  �       o   �� ���        ������  ����������������        ��� ��    x                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    x                    ����    �  �       o   �� ���        ������  ����������������        ��� ��    <                    ����    �  �       p   �� ���        ������  ����������������        ��� ��    <  
                  ����    �  �       p   �� ���        ������  ����������������        ��� ��    <                    ����    �  �        p   �� ���        ������  ����������������        ��� ��    <                    ����    �  �     !  p   �� ���        ������  ����������������        ��� ��    x                    ����    �  �     "  p   �� ���        ������  ����������������        ��� ��    x  
                  ����    �  �     #  p   �� ���        ������  ����������������        ��� ��    x                    ����    �  �     $  p   �� ���        ������  ����������������        ��� ��    x                    ����    �  �     %  p   �� ���        ������  ����������������        ��� ��'                        ����    �  �     &  q   �� ���        ������  ����������������        ��� ��(                        ����    �  �     '  r   �� ���        ������  ����������������        ��� ��                           ����    �  �     (  s   �� ���        ������  ����������������        ��� ��         
                  ����    �  �     )  s   �� ���        ������  ����������������        ��� ��                           ����    �  �     *  s   �� ���        ������  ����������������        ��� ��                           ����    �  �     +  s   �� ���        ������  ����������������        ��� ��                           ����    �  �     ,  t   �� ���        ������  ����������������        ��� ��         
                  ����    �  �     -  t   �� ���        ������  ����������������        ��� ��                           ����    �  �     .  t   �� ���        ������  ����������������        ��� ��                           ����    �  �     /  t   �� ���        ������  ����������������        ��� ��                         ����    �  �     0  u   �� ���        ������  ����������������        ��� ��       
                  ����    �  �     1  u   �� ���        ������  ����������������        ��� ��                         ����    �  �     2  u   �� ���        ������  ����������������        ��� ��                         ����    �  �     3  u   �� ���        ������  ����������������        ��� ��                         ����    �  �     4  u   �� ���        ������  ����������������        ��� ��       
                  ����    �  �     5  u   �� ���        ������  ����������������        ��� ��                         ����    �  �     6  u   �� ���        ������  ����������������        ��� ��                         ����    �  �     7  u   �� ���        ������  ����������������        ��� ��                        ����    �  �     8  v   �� ���        ������  ����������������        ��� ��      
                  ����    �  �     9  v   �� ���        ������  ����������������        ��� ��                        ����    �  �     :  v   �� ���        ������  ����������������        ��� ��                        ����    �  �     ;  v   �� ���        ������  ����������������        ��� ��                        ����    �  �     <  v   �� ���        ������  ����������������        ��� ��      
                  ����    �  �     =  v   �� ���        ������  ����������������        ��� ��                        ����    �  �     >  v   �� ���        ������  ����������������        ��� ��                        ����    �  �     ?  v   �� ���        ������  ����������������        ��� ��d P                        ����    �  �     @  w   �� ���        ������  ����������������        ��� ��d P      
                  ����    �  �     A  w   �� ���        ������  ����������������        ��� ��d P                        ����    �  �     B  w   �� ���        ������  ����������������        ��� ��d P                        ����    �  �     C  w   �� ���        ������  ����������������        ��� ��                             �5w    �  �     D      �� ���        ������  ����������������        ��� ��                            ����    �  �     E  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     F  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     G  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     H  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     I  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     J  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     K  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     L  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     M  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     N  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     O  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     P  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     Q  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     R  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     S  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     T  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     U  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     V  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     W  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     X  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     Y  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     Z  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     [  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     \  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     ]  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     ^  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     _  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     `  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     a  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     b  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     c  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     d  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     e  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     f  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     g  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     h  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     i  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     j  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     k  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     l  �   �� ���        ������  ����������������        ��� ��)                       ����    �  �     m  x   �� ���        ������  ����������������        ��� ��)                       ����    �  �     n  x   �� ���        ������  ����������������        ��� ��)     
                  ����    �  �     o  x   �� ���        ������  ����������������        ��� ��*                        ����    �  �     p  y   �� ���        ������  ����������������        ��� ��*                        ����    �  �     q  y   �� ���        ������  ����������������        ��� ��*      
                  ����    �  �     r  y   �� ���        ������  ����������������        ��� ��                          ����    �  �     s  w   �� ���        ������  ����������������        ��� ��        7                  ����    �  �     t  w   �� ���        ������  ����������������        ��� ��        x                  ����    �  �     u  w   �� ���        ������  ����������������        ��� ��        �                  ����    �  �     v  w   �� ���        ������  ����������������          ����[2    d                 �  �                   M    �������c   ������������b            ���$�]2    i                 �  �                  M    �������c   ������������b            ���)�_2    n                 :  �                  M    �������c   ������������b            ���.�a2    s                 �  �                  M   �������c   ������������b            ���3�c2    x                 �  �                  M   �������c   ������������b            ���8�e2    }                 H   !                  M   �������c   ������������b            ���=�g2    �                 �  �"                  M   �������c   ������������b            ���B�i2    �                 �  �#                  M   �������c   ������������b            ���G�k2    �                 V	  X%                  M   �������c   ������������b            ���L�m2    �                 �	  �&         	         M   �������c   ������������b            ���[�2        d             �  �e        p       h   N    �������c   ������������c            ���]�$2        i             �  <i        p      h   N    �������c   ������������c            ���_�)2        n                �l        p      h   N    �������c   ������������c            ���a�.2        s             �  Dp        p      h   N   �������c   ������������c            ���c�32        x             L  �s        p      h   N   �������c   ������������c            ���e�82        }             �  Lw        p      h   N   �������c   ������������c            ���g�=2        �             x  �z        p      h   N   �������c   ������������c            ���i�B2        �               T~        p      h   N   �������c   ������������c            ���k�G2        �             �  ؁        p      h   N   �������c   ������������c            ���m�L2        �             :  \�        p 	     h   N   �������c   ������������c             ��
2      K K             �  �9        �       �   O    �������c   ������������d             ��
2      M O               (<        �      �   O    �������c   ������������d             �	�	
2      O S             �  �>        �      �   O    �������c   ������������d             ��
2      Q W             �  �@        �      �   O   �������c   ������������d             ��
2      S [             p  0C        �      �   O   �������c   ������������d             ��
2      U _             �  �E        �      �   O   �������c   ������������d             ��
2      W c             `  �G        �      �   O   �������c   ������������d             ��
2      Y g             �  8J        �      �   O   �������c   ������������d             �!�!
2      [ k             P  �L        �      �   O   �������c   ������������d             �%�%
2      ] o             �  �N        � 	     �   O   �������c   ������������d             ��=2    K K               v  �        �       �   �    �������c   ������������e             ��?2    M N               �  @        �      �   �    �������c   ������������e             ��A2    O Q               *  �         �      �   �    �������c   ������������e             ��C2    Q T               �  "        �      �   �   �������c   ������������e             ��E2    S W               �  x#        �      �   �   �������c   ������������e             $��G2    U Z               8	  �$        �      �   �   �������c   ������������e             )��I2    W ]               �	  H&        �      �   �   �������c   ������������e             .��K2    Y `               �	  �'        �      �   �   �������c   ������������e             3��M2    [ c               F
  )        �      �   �   �������c   ������������e             8��O2    ] f               �
  �*        � 	     �   �   �������c   ������������e            ���/�/2    ,d d 2           �  "        A       >       �������c   ������������f            ���J�J2    1i i 7           �  �        A      >       �������c   ������������f            ���e�e2    6n n <           .  �        A      >       �������c   ������������f            ������2    ;s s A           j  >        A      >      �������c   ������������f            ������2    @x x F           �  �        A      >      �������c   ������������f            ����2    E} } K           �  �        A      >      �������c   ������������f            ��)�)�2    J� � P             Z        A      >      �������c   ������������f            ��C�C�2    O� � U           Z          A      >      �������c   ������������f            ��]]2    T� � Z           �  �        A      >      �������c   ������������f            ��w"w"2    Y� � _           �  v        A 	     >      �������c   ������������f            �����2    ,d d 2           .  �        W       S       �������c   ������������g            ��'��2    1i i 7           j  >        W      S       �������c   ������������g            ��C�+�2    6n n <           �  �        W      S       �������c   ������������g            ��_C�2    ;s s A           �  �        W      S      �������c   ������������g            ��{![�2    @x x F             Z        W      S      �������c   ������������g            ���>s2    E} } K           Z          W      S      �������c   ������������g            ���[�12    J� � P           �  �        W      S      �������c   ������������g            ���x�K2    O� � U           �  v        W      S      �������c   ������������g            �����e2    T� � Z             *        W      S      �������c   ������������g            ����2    Y� � _           J  �        W 	     S      �������c   ������������g            ���/�T2    d d ,2           �  ��        q       k       �������c   ������������h            ���G�s2    i i 17           F  �        q      k       �������c   ������������h            ���_��2    n n 6<           �  ֵ        q      k       �������c   ������������h            ���w�2    s s ;A           �  º        q      k      �������c   ������������h            ����3�2    x x @F           b  ��        q      k      �������c   ������������h            ����Q�2    } } EK             ��        q      k      �������c   ������������h            ���o2    � � JP           �  ��        q      k      �������c   ������������h            ��#��-2    � � OU           ~  r�        q      k      �������c   ������������h            ��:��L2    � � TZ           2  ^�        q      k      �������c   ������������h            ��Q�k2    � � Y_           �  J�        q 	     k      �������c   ������������h             S�S�
2    ,d d 2           �  �i        �       �       �������c   ������������i             l
l

2    1i i 7           >  tm        �      �       �������c   ������������i             �%�%
2    6n n <           �  �p        �      �       �������c   ������������i             �@�@
2    ;s s A           j  |t        �      �      �������c   ������������i             �[�[
2    @x x F               x        �      �      �������c   ������������i             �v�v
2    E} } K           �  �{        �      �      �������c   ������������i             ����
2    J� � P           ,          �      �      �������c   ������������i             ��
2    O� � U           �  ��        �      �      �������c   ������������i             ��
2    T� � Z           X  �        �      �      �������c   ������������i             4�4�
2    Y� � _           �  ��        � 	     �      �������c   ������������i             a�/2    d ,d 2             (<        �       �       �������c   ������������j             ~6�G2    i 1i 7           �  �>        �      �       �������c   ������������j             �T�_2    n 6n <           �  �@        �      �       �������c   ������������j             �r�w2    s ;s A           p  0C        �      �      �������c   ������������j             ����2    x @x F           �  �E        �      �      �������c   ������������j             ����2    } E} K           `  �G        �      �      �������c   ������������j             ��2    � J� P           �  8J        �      �      �������c   ������������j             ,�#�2    � O� U           P  �L        �      �      �������c   ������������j             I:�2    � T� Z           �  �N        �      �      �������c   ������������j             f&Q2    � Y� _           @  @Q        � 	     �      �������c   ������������j         ����   / 0          � d               \  (n        )        ��        ����c   ������������k         ����   2 3          � g               �  �q        )       ��        ����c   ������������k         ����   5 6          � j               �  0u        )       ��        ����c   ������������k         ����   8 9          � m                 �x        )       ��       ����c   ������������k         ����   ; <          � p               �  8|        )       ��       ����c   ������������k         ����   > ?          � s               J  �        )       ��       ����c   ������������k         ����   A B          � v               �  @�        )       ��       ����c   ������������k         ����   D E          � y               v  Ć        )       ��       ����c   ������������k         ����   G H          � |                 H�        )       ��       ����c   ������������k         ����   J K          �                �  ̍        )	       ��       ����c   ������������k         ����  - .          � d               �          �        ��        ����c   ������������l         ����  0 1          � g               �  �        �       ��        ����c   ������������l         ����  3 4          � j               *  ~	        �       ��        ����c   ������������l         ����  6 7          � m               f  2
        �       ��       ����c   ������������l         ����  9 :          � p               �  �
        �       ��       ����c   ������������l         ����  < =          � s               �  �        �       ��       ����c   ������������l         ����  ? @          � v                 N        �       ��       ����c   ������������l         ����  B C          � y               V          �       ��       ����c   ������������l         ����  E F          � |               �  �        �       ��       ����c   ������������l         ����  H I          �                �  j        �	       ��       ����c   ������������l         ����  . /          � d               N  �                 ��        ����c   ������������m         ����  1 2          � g               �  �                ��        ����c   ������������m         ����  4 5          � j               �  R                ��        ����c   ������������m         ����  7 8          � m                 	                ��       ����c   ������������m         ����  : ;          � p               >  �	                ��       ����c   ������������m         ����  = >          � s               z  n
                ��       ����c   ������������m         ����  @ A          � v               �  "                ��       ����c   ������������m         ����  C D          � y               �  �                ��       ����c   ������������m         ����  F G          � |               .  �                ��       ����c   ������������m         ����  I J          �                j  >         	       ��       ����c   ������������m         ����  - .          � d               V	          f        ��        ����c   ������������n         ����  0 1          � g               �	  �        f       ��        ����c   ������������n         ����  3 4          � j               �	  j        f       ��        ����c   ������������n         ����  6 7          � m               

          f       ��       ����c   ������������n         ����  9 :          � p               F
  �        f       ��       ����c   ������������n         ����  < =          � s               �
  �        f       ��       ����c   ������������n         ����  ? @          � v               �
  :         f       ��       ����c   ������������n         ����  B C          � y               �
  �         f       ��       ����c   ������������n         ����  E F          � |               6  �!        f       ��       ����c   ������������n         ����  H I          �                r  V"        f	       ��       ����c   ������������n         ����  0 1          � d               �  R        �        ��        ����c   ������������o         ����  3 4          � g                         �       ��        ����c   ������������o         ����  6 7          � j               >  �        �       ��        ����c   ������������o         ����  9 :          � m               z  n        �       ��       ����c   ������������o         ����  < =          � p               �  "        �       ��       ����c   ������������o         ����  ? @          � s               �  �        �       ��       ����c   ������������o         ����  B C          � v               .	  �        �       ��       ����c   ������������o         ����  E F          � y               j	  >        �       ��       ����c   ������������o         ����  H I          � |               �	  �        �       ��       ����c   ������������o         ����  K L          �                �	  �        �	       ��       ����c   ������������o         ����  . /          � d               6  �        2        ��         ����c   ������������p         ����  1 2          � g               r  V        2       ��         ����c   ������������p         ����  4 5          � j               �  
        2       ��         ����c   ������������p         ����  7 8          � m               �  �        2       ��        ����c   ������������p         ����  : ;          � p               &  r        2       ��        ����c   ������������p         ����  = >          � s               b  &        2       ��        ����c   ������������p         ����  @ A          � v               �  �        2       ��        ����c   ������������p         ����  C D          � y               �  �        2       ��        ����c   ������������p         ����  F G          � |                 B        2       ��        ����c   ������������p         ����  I J          �                R  �        2	       ��        ����c   ������������p         ����  / 0          � d               �
  �         �      �   �        ����c   ������������q         ����  2 3          � g               "  f!        �     �   �        ����c   ������������q         ����  5 6          � j               ^  "        �     �   �        ����c   ������������q         ����  8 9          � m               �  �"        �     �   �       ����c   ������������q         ����  ; <          � p               �  �#        �     �   �       ����c   ������������q         ����  > ?          � s                 6$        �     �   �       ����c   ������������q         ����  A B          � v               N  �$        �     �   �       ����c   ������������q         ����  D E          � y               �  �%        �     �   �       ����c   ������������q         ����  G H          � |               �  R&        �     �   �       ����c   ������������q         ����  J K          �                  '        �	     �   �       ����c   ������������q         ����   % &            d �             \  (n        =        ��        ����c   ������������r         ����   ( )            g �             �  �q        =       ��        ����c   ������������r         ����   + ,            j �             �  0u        =       ��        ����c   ������������r         ����   . /            m �               �x        =       ��       ����c   ������������r         ����   1 2            p �             �  8|        =       ��       ����c   ������������r         ����   4 5            s �             J  �        =       ��       ����c   ������������r         ����   7 8            v �             �  @�        =       ��       ����c   ������������r         ����   : ;            y �             v  Ć        =       ��       ����c   ������������r         ����   = >            | �               H�        =       ��       ����c   ������������r         ����   @ A             �             �  ̍        =	       ��       ����c   ������������r         ����  $ %            d �             �          �        ��
        ����c   ������������s         ����  ' (            g �             �  �        �       ��
        ����c   ������������s         ����  * +            j �             *  ~	        �       ��
        ����c   ������������s         ����  - .            m �             f  2
        �       ��
       ����c   ������������s         ����  0 1            p �             �  �
        �       ��
       ����c   ������������s         ����  3 4            s �             �  �        �       ��
       ����c   ������������s         ����  6 7            v �               N        �       ��
       ����c   ������������s         ����  9 :            y �             V          �       ��
       ����c   ������������s         ����  < =            | �             �  �        �       ��
       ����c   ������������s         ����  ? @             �             �  j        �	       ��
       ����c   ������������s         ����  $ %            d �             N  �                ��        ����c   ������������t         ����  ' (            g �             �  �               ��        ����c   ������������t         ����  * +            j �             �  R               ��        ����c   ������������t         ����  - .            m �               	               ��       ����c   ������������t         ����  0 1            p �             >  �	               ��       ����c   ������������t         ����  3 4            s �             z  n
               ��       ����c   ������������t         ����  6 7            v �             �  "               ��       ����c   ������������t         ����  9 :            y �             �  �               ��       ����c   ������������t         ����  < =            | �             .  �               ��       ����c   ������������t         ����  ? @             �             j  >        	       ��       ����c   ������������t         ����  $ %            d �             V	          w        ��        ����c   ������������u         ����  ' (            g �             �	  �        w       ��        ����c   ������������u         ����  * +            j �             �	  j        w       ��        ����c   ������������u         ����  - .            m �             

          w       ��       ����c   ������������u         ����  0 1            p �             F
  �        w       ��       ����c   ������������u         ����  3 4            s �             �
  �        w       ��       ����c   ������������u         ����  6 7            v �             �
  :         w       ��       ����c   ������������u         ����  9 :            y �             �
  �         w       ��       ����c   ������������u         ����  < =            | �             6  �!        w       ��       ����c   ������������u         ����  ? @             �             r  V"        w	       ��       ����c   ������������u         ����  % &            d �             �  R        �        ��        ����c   ������������v         ����  ( )            g �                       �       ��        ����c   ������������v         ����  + ,            j �             >  �        �       ��        ����c   ������������v         ����  . /            m �             z  n        �       ��       ����c   ������������v         ����  1 2            p �             �  "        �       ��       ����c   ������������v         ����  4 5            s �             �  �        �       ��       ����c   ������������v         ����  7 8            v �             .	  �        �       ��       ����c   ������������v         ����  : ;            y �             j	  >        �       ��       ����c   ������������v         ����  = >            | �             �	  �        �       ��       ����c   ������������v         ����  @ A             �             �	  �        �	       ��       ����c   ������������v         ����  $ %            d �             6  �        C        ��"        ����c   ������������w         ����  ' (            g �             r  V        C       ��"        ����c   ������������w         ����  * +            j �             �  
        C       ��"        ����c   ������������w         ����  - .            m �             �  �        C       ��"       ����c   ������������w         ����  0 1            p �             &  r        C       ��"       ����c   ������������w         ����  3 4            s �             b  &        C       ��"       ����c   ������������w         ����  6 7            v �             �  �        C       ��"       ����c   ������������w         ����  9 :            y �             �  �        C       ��"       ����c   ������������w         ����  < =            | �               B        C       ��"       ����c   ������������w         ����  ? @             �             R  �        C	       ��"       ����c   ������������w         ����  % &            d �             �
  �         �      �   �        ����c   ������������x         ����  ( )            g �             "  f!        �     �   �        ����c   ������������x         ����  + ,            j �             ^  "        �     �   �        ����c   ������������x         ����  . /            m �             �  �"        �     �   �       ����c   ������������x         ����  1 2            p �             �  �#        �     �   �       ����c   ������������x         ����  4 5            s �               6$        �     �   �       ����c   ������������x         ����  7 8            v �             N  �$        �     �   �       ����c   ������������x         ����  : ;            y �             �  �%        �     �   �       ����c   ������������x         ����  = >            | �             �  R&        �     �   �       ����c   ������������x         ����  @ A             �               '        �	     �   �       ����c   ������������x         ����   $ %          �   �             \  (n        Q        ��        ����c   ������������y         ����   ' (          �   �             �  �q        Q       ��        ����c   ������������y         ����   * +          �   �             �  0u        Q       ��        ����c   ������������y         ����   - .          �   �               �x        Q       ��       ����c   ������������y         ����   0 1          �   �             �  8|        Q       ��       ����c   ������������y         ����   3 4          �   �             J  �        Q       ��       ����c   ������������y         ����   6 7          �   �             �  @�        Q       ��       ����c   ������������y         ����   9 :          �   �             v  Ć        Q       ��       ����c   ������������y         ����   < =          �   �               H�        Q       ��       ����c   ������������y         ����   ? @          �   �             �  ̍        Q	       ��       ����c   ������������y         ����  # $          �   �             �          �        ��        ����c   ������������z         ����  & '          �   �             �  �        �       ��        ����c   ������������z         ����  ) *          �   �             *  ~	        �       ��        ����c   ������������z         ����  , -          �   �             f  2
        �       ��       ����c   ������������z         ����  / 0          �   �             �  �
        �       ��       ����c   ������������z         ����  2 3          �   �             �  �        �       ��       ����c   ������������z         ����  5 6          �   �               N        �       ��       ����c   ������������z         ����  8 9          �   �             V          �       ��       ����c   ������������z         ����  ; <          �   �             �  �        �       ��       ����c   ������������z         ����  > ?          �   �             �  j        �	       ��       ����c   ������������z         ����  # $          �   �             N  �        "        ��        ����c   ������������{         ����  & '          �   �             �  �        "       ��        ����c   ������������{         ����  ) *          �   �             �  R        "       ��        ����c   ������������{         ����  , -          �   �               	        "       ��       ����c   ������������{         ����  / 0          �   �             >  �	        "       ��       ����c   ������������{         ����  2 3          �   �             z  n
        "       ��       ����c   ������������{         ����  5 6          �   �             �  "        "       ��       ����c   ������������{         ����  8 9          �   �             �  �        "       ��       ����c   ������������{         ����  ; <          �   �             .  �        "       ��       ����c   ������������{         ����  > ?          �   �             j  >        "	       ��       ����c   ������������{         ����  # $          �   �             V	          �        ��        ����c   ������������|         ����  & '          �   �             �	  �        �       ��        ����c   ������������|         ����  ) *          �   �             �	  j        �       ��        ����c   ������������|         ����  , -          �   �             

          �       ��       ����c   ������������|         ����  / 0          �   �             F
  �        �       ��       ����c   ������������|         ����  2 3          �   �             �
  �        �       ��       ����c   ������������|         ����  5 6          �   �             �
  :         �       ��       ����c   ������������|         ����  8 9          �   �             �
  �         �       ��       ����c   ������������|         ����  ; <          �   �             6  �!        �       ��       ����c   ������������|         ����  > ?          �   �             r  V"        �	       ��       ����c   ������������|         ����  $ %          �   �             �  R        �        ��        ����c   ������������}         ����  ' (          �   �                       �       ��        ����c   ������������}         ����  * +          �   �             >  �        �       ��        ����c   ������������}         ����  - .          �   �             z  n        �       ��       ����c   ������������}         ����  0 1          �   �             �  "        �       ��       ����c   ������������}         ����  3 4          �   �             �  �        �       ��       ����c   ������������}         ����  6 7          �   �             .	  �        �       ��       ����c   ������������}         ����  9 :          �   �             j	  >        �       ��       ����c   ������������}         ����  < =          �   �             �	  �        �       ��       ����c   ������������}         ����  ? @          �   �             �	  �        �	       ��       ����c   ������������}         ����  # $          �   �             6  �        T        ��$        ����c   ������������~         ����  & '          �   �             r  V        T       ��$        ����c   ������������~         ����  ) *          �   �             �  
        T       ��$        ����c   ������������~         ����  , -          �   �             �  �        T       ��$       ����c   ������������~         ����  / 0          �   �             &  r        T       ��$       ����c   ������������~         ����  2 3          �   �             b  &        T       ��$       ����c   ������������~         ����  5 6          �   �             �  �        T       ��$       ����c   ������������~         ����  8 9          �   �             �  �        T       ��$       ����c   ������������~         ����  ; <          �   �               B        T       ��$       ����c   ������������~         ����  > ?          �   �             R  �        T	       ��$       ����c   ������������~         ����  $ %          �   �             �
  �         �      �   �        ����c   ������������         ����  ' (          �   �             "  f!        �     �   �        ����c   ������������         ����  * +          �   �             ^  "        �     �   �        ����c   ������������         ����  - .          �   �             �  �"        �     �   �       ����c   ������������         ����  0 1          �   �             �  �#        �     �   �       ����c   ������������         ����  3 4          �   �               6$        �     �   �       ����c   ������������         ����  6 7          �   �             N  �$        �     �   �       ����c   ������������         ����  9 :          �   �             �  �%        �     �   �       ����c   ������������         ����  < =          �   �             �  R&        �     �   �       ����c   ������������         ����  ? @          �   �               '        �	     �   �       ����c   ������������         ����                d �             \  (n        e        ���        ����c   �������������         ����                 g �             �  �q        e       ���        ����c   �������������         ����   " #            j �             �  0u        e       ���        ����c   �������������         ����   % &            m �               �x        e       ���       ����c   �������������         ����   ( )            p �             �  8|        e       ���       ����c   �������������         ����   + ,            s �             J  �        e       ���       ����c   �������������         ����   . /            v �             �  @�        e       ���       ����c   �������������         ����   1 2            y �             v  Ć        e       ���       ����c   �������������         ����   4 5            | �               H�        e       ���       ����c   �������������         ����   7 8             �             �  ̍        e	       ���       ����c   �������������         ����               d �             �          �        ���        ����c   �������������         ����               g �             �  �        �       ���        ����c   �������������         ����  ! "            j �             *  ~	        �       ���        ����c   �������������         ����  $ %            m �             f  2
        �       ���       ����c   �������������         ����  ' (            p �             �  �
        �       ���       ����c   �������������         ����  * +            s �             �  �        �       ���       ����c   �������������         ����  - .            v �               N        �       ���       ����c   �������������         ����  0 1            y �             V          �       ���       ����c   �������������         ����  3 4            | �             �  �        �       ���       ����c   �������������         ����  6 7             �             �  j        �	       ���       ����c   �������������         ����               d �             N  �        3        ���        ����c   �������������         ����               g �             �  �        3       ���        ����c   �������������         ����  ! "            j �             �  R        3       ���        ����c   �������������         ����  $ %            m �               	        3       ���       ����c   �������������         ����  ' (            p �             >  �	        3       ���       ����c   �������������         ����  * +            s �             z  n
        3       ���       ����c   �������������         ����  - .            v �             �  "        3       ���       ����c   �������������         ����  0 1            y �             �  �        3       ���       ����c   �������������         ����  3 4            | �             .  �        3       ���       ����c   �������������         ����  6 7             �             j  >        3	       ���       ����c   �������������         ����               d �             V	          �        ���        ����c   �������������         ����               g �             �	  �        �       ���        ����c   �������������         ����  ! "            j �             �	  j        �       ���        ����c   �������������         ����  $ %            m �             

          �       ���       ����c   �������������         ����  ' (            p �             F
  �        �       ���       ����c   �������������         ����  * +            s �             �
  �        �       ���       ����c   �������������         ����  - .            v �             �
  :         �       ���       ����c   �������������         ����  0 1            y �             �
  �         �       ���       ����c   �������������         ����  3 4            | �             6  �!        �       ���       ����c   �������������         ����  6 7             �             r  V"        �	       ���       ����c   �������������         ����               d �             �  R        �        ���        ����c   �������������         ����                g �                       �       ���        ����c   �������������         ����  " #            j �             >  �        �       ���        ����c   �������������         ����  % &            m �             z  n        �       ���       ����c   �������������         ����  ( )            p �             �  "        �       ���       ����c   �������������         ����  + ,            s �             �  �        �       ���       ����c   �������������         ����  . /            v �             .	  �        �       ���       ����c   �������������         ����  1 2            y �             j	  >        �       ���       ����c   �������������         ����  4 5            | �             �	  �        �       ���       ����c   �������������         ����  7 8             �             �	  �        �	       ���       ����c   �������������         ����               d �             6  �        e        ���        ����c   �������������         ����               g �             r  V        e       ���        ����c   �������������         ����  ! "            j �             �  
        e       ���        ����c   �������������         ����  $ %            m �             �  �        e       ���       ����c   �������������         ����  ' (            p �             &  r        e       ���       ����c   �������������         ����  * +            s �             b  &        e       ���       ����c   �������������         ����  - .            v �             �  �        e       ���       ����c   �������������         ����  0 1            y �             �  �        e       ���       ����c   �������������         ����  3 4            | �               B        e       ���       ����c   �������������         ����  6 7             �             R  �        e	       ���       ����c   �������������         ����               d �             �
  �         �      �   |        ����c   �������������         ����    !            g �             "  f!        �     �   |        ����c   �������������         ����  # $            j �             ^  "        �     �   |        ����c   �������������         ����  & '            m �             �  �"        �     �   |       ����c   �������������         ����  ) *            p �             �  �#        �     �   |       ����c   �������������         ����  , -            s �               6$        �     �   |       ����c   �������������         ����  / 0            v �             N  �$        �     �   |       ����c   �������������         ����  2 3            y �             �  �%        �     �   |       ����c   �������������         ����  5 6            | �             �  R&        �     �   |       ����c   �������������         ����  8 9             �               '        �	     �   |       ����c   �������������         ����   % &          d �               �  �        w        ���        ����c   �������������         ����   ( )          g �                 0         w       ���        ����c   �������������         ����   + ,          j �               f  �!        w       ���        ����c   �������������         ����   . /          m �               �   #        w       ���       ����c   �������������         ����   1 2          p �               	  h$        w       ���       ����c   �������������         ����   4 5          s �               t	  �%        w       ���       ����c   �������������         ����   7 8          v �               �	  8'        w       ���       ����c   �������������         ����   : ;          y �               (
  �(        w       ���       ����c   �������������         ����   = >          | �               �
  *        w       ���       ����c   �������������         ����   @ A           �               �
  p+        w	       ���       ����c   �������������         ����  $ %          d �               N  �        D        ���        ����c   �������������         ����  ' (          g �               �  �        D       ���        ����c   �������������         ����  * +          j �               �  R        D       ���        ����c   �������������         ����  - .          m �                 	        D       ���       ����c   �������������         ����  0 1          p �               >  �	        D       ���       ����c   �������������         ����  3 4          s �               z  n
        D       ���       ����c   �������������         ����  6 7          v �               �  "        D       ���       ����c   �������������         ����  9 :          y �               �  �        D       ���       ����c   �������������         ����  < =          | �               .  �        D       ���       ����c   �������������         ����  ? @           �               j  >        D	       ���       ����c   �������������         ����  $ %          d �               �          �        ���        ����c   �������������         ����  ' (          g �               �  �        �       ���        ����c   �������������         ����  * +          j �               *  ~	        �       ���        ����c   �������������         ����  - .          m �               f  2
        �       ���       ����c   �������������         ����  0 1          p �               �  �
        �       ���       ����c   �������������         ����  3 4          s �               �  �        �       ���       ����c   �������������         ����  6 7          v �                 N        �       ���       ����c   �������������         ����  9 :          y �               V          �       ���       ����c   �������������         ����  < =          | �               �  �        �       ���       ����c   �������������         ����  ? @           �               �  j        �	       ���       ����c   �������������         ����  $ %          d �               V	          �        ���        ����c   �������������         ����  ' (          g �               �	  �        �       ���        ����c   �������������         ����  * +          j �               �	  j        �       ���        ����c   �������������         ����  - .          m �               

          �       ���       ����c   �������������         ����  0 1          p �               F
  �        �       ���       ����c   �������������         ����  3 4          s �               �
  �        �       ���       ����c   �������������         ����  6 7          v �               �
  :         �       ���       ����c   �������������         ����  9 :          y �               �
  �         �       ���       ����c   �������������         ����  < =          | �               6  �!        �       ���       ����c   �������������         ����  ? @           �               r  V"        �	       ���       ����c   �������������         ����  $ %          d �               6  �        v        ���        ����c   �������������         ����  ' (          g �               r  V        v       ���        ����c   �������������         ����  * +          j �               �  
        v       ���        ����c   �������������         ����  - .          m �               �  �        v       ���       ����c   �������������         ����  0 1          p �               &  r        v       ���       ����c   �������������         ����  3 4          s �               b  &        v       ���       ����c   �������������         ����  6 7          v �               �  �        v       ���       ����c   �������������         ����  9 :          y �               �  �        v       ���       ����c   �������������         ����  < =          | �                 B        v       ���       ����c   �������������         ����  ? @           �               R  �        v	       ���       ����c   �������������         ����  % &          d �               �  R                ���        ����c   �������������         ����  ( )          g �                                ���        ����c   �������������         ����  + ,          j �               >  �               ���        ����c   �������������         ����  . /          m �               z  n               ���       ����c   �������������         ����  1 2          p �               �  "               ���       ����c   �������������         ����  4 5          s �               �  �               ���       ����c   �������������         ����  7 8          v �               .	  �               ���       ����c   �������������         ����  : ;          y �               j	  >               ���       ����c   �������������         ����  = >          | �               �	  �               ���       ����c   �������������         ����  @ A           �               �	  �        	       ���       ����c   �������������         ����    $ %            � �             �  �        �        ��         ����c   �������������         ����    ' (            � �               0         �       ��         ����c   �������������         ����    * +            � �             f  �!        �       ��         ����c   �������������         ����    - .            � �             �   #        �       ��        ����c   �������������         ����    0 1            � �             	  h$        �       ��        ����c   �������������         ����    3 4            � �             t	  �%        �       ��        ����c   �������������         ����    6 7            � �             �	  8'        �       ��        ����c   �������������         ����    9 :            � �             (
  �(        �       ��        ����c   �������������         ����    < =            � �             �
  *        �       ��        ����c   �������������         ����    ? @            � �             �
  p+        �	       ��        ����c   �������������         ����   # $            � �             �          �        ��        ����c   �������������         ����   & '            � �             �  �        �       ��        ����c   �������������         ����   ) *            � �             *  ~	        �       ��        ����c   �������������         ����   , -            � �             f  2
        �       ��       ����c   �������������         ����   / 0            � �             �  �
        �       ��       ����c   �������������         ����   2 3            � �             �  �        �       ��       ����c   �������������         ����   5 6            � �               N        �       ��       ����c   �������������         ����   8 9            � �             V          �       ��       ����c   �������������         ����   ; <            � �             �  �        �       ��       ����c   �������������         ����   > ?            � �             �  j        �	       ��       ����c   �������������         ����   # $            � �             N  �        U        ��        ����c   �������������         ����   & '            � �             �  �        U       ��        ����c   �������������         ����   ) *            � �             �  R        U       ��        ����c   �������������         ����   , -            � �               	        U       ��       ����c   �������������         ����   / 0            � �             >  �	        U       ��       ����c   �������������         ����   2 3            � �             z  n
        U       ��       ����c   �������������         ����   5 6            � �             �  "        U       ��       ����c   �������������         ����   8 9            � �             �  �        U       ��       ����c   �������������         ����   ; <            � �             .  �        U       ��       ����c   �������������         ����   > ?            � �             j  >        U	       ��       ����c   �������������         ����   # $            � �             V	          �        ��        ����c   �������������         ����   & '            � �             �	  �        �       ��        ����c   �������������         ����   ) *            � �             �	  j        �       ��        ����c   �������������         ����   , -            � �             

          �       ��       ����c   �������������         ����   / 0            � �             F
  �        �       ��       ����c   �������������         ����   2 3            � �             �
  �        �       ��       ����c   �������������         ����   5 6            � �             �
  :         �       ��       ����c   �������������         ����   8 9            � �             �
  �         �       ��       ����c   �������������         ����   ; <            � �             6  �!        �       ��       ����c   �������������         ����   > ?            � �             r  V"        �	       ��       ����c   �������������         ����   $ %            � �             �  R        !        ��        ����c   �������������         ����   ' (            � �                       !       ��        ����c   �������������         ����   * +            � �             >  �        !       ��        ����c   �������������         ����   - .            � �             z  n        !       ��       ����c   �������������         ����   0 1            � �             �  "        !       ��       ����c   �������������         ����   3 4            � �             �  �        !       ��       ����c   �������������         ����   6 7            � �             .	  �        !       ��       ����c   �������������         ����   9 :            � �             j	  >        !       ��       ����c   �������������         ����   < =            � �             �	  �        !       ��       ����c   �������������         ����   ? @            � �             �	  �        !	       ��       ����c   �������������         ����   # $            � �             6  �        �        ��        ����c   �������������         ����   & '            � �             r  �        �       ��        ����c   �������������         ����   ) *            � �             �  �        �       ��        ����c   �������������         ����   , -            � �             �  �        �       ��       ����c   �������������         ����   / 0            � �             &  �        �       ��       ����c   �������������         ����   2 3            � �             b  �        �       ��       ����c   �������������         ����   5 6            � �             �  �        �       ��       ����c   �������������         ����   8 9            � �             �  �        �       ��       ����c   �������������         ����   ; <            � �               �        �       ��       ����c   �������������         ����   > ?            � �             R  �        �	       ��       ����c   �������������         ����   $ %            � �             �
  �        �      �           ����c   �������������         ����   ' (            � �             "  �        �     �           ����c   �������������         ����   * +            � �             ^  �        �     �           ����c   �������������         ����   - .            � �             �  �        �     �          ����c   �������������         ����   0 1            � �             �  �        �     �          ����c   �������������         ����   3 4            � �               �        �     �          ����c   �������������         ����   6 7            � �             N  �        �     �          ����c   �������������         ����   9 :            � �             �  �        �     �          ����c   �������������         ����   < =            � �             �  �        �     �          ����c   �������������         ����   ? @            � �               �        �	     �          ����c   �������������          ��� ��                       ����    �  �     w  z   �� ���        ������  ����������������        ��� �� (                      ����    �  �     x  z   �� ���        ������  ����������������        ��� ��                       ����    �  �     y  {   �� ���        ������  ����������������        ��� �� (                      ����    �  �     z  {   �� ���        ������  ����������������        ��� ��                       ����    �  �     {  |   �� ���        ������  ����������������        ��� �� (                      ����    �  �     |  |   �� ���        ������  ����������������        ��� ��                       ����    �  �     }  }   �� ���        ������  ����������������        ��� �� (                      ����    �  �     ~  }   �� ���        ������  ����������������       ����                               ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                                ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                              ����                         ��        ����c   �������������         ����                               ����                         ��        ����c   �������������          ��d ��                         �   L  �  �          ��. ��<        ������  ����������������        ��d ��                         �   �  �  �     �     ��. ��=        ������  ����������������        ��d ��  (        
               �   8  �  �     �     ��. ��>        ������  ����������������        ��d ��  2                       �   �  �  �     �     ��. ��?        ������  ����������������        ��d ��  P        &               �   P�  �  �     �     ��. ��#        ������  ����������������        ��d ��  d        <               �   �$ �  �     �     ��. ��$        ������  ����������������        ��e ��                         �   L  �  �     �     ��/ ��@        ������  ����������������        ��e ��                         �   �  �  �     �     ��/ ��A        ������  ����������������        ��e ��  (        
               �   8  �  �     �     ��/ ��B        ������  ����������������        ��e ��  2                       �   �  �  �     �     ��/ ��C        ������  ����������������        ��e ��  P        &               �   P�  �  �     �     ��/ ��%        ������  ����������������        ��e ��  d        <               �   �$ �  �     �     ��/ ��&        ������  ����������������        ��d ��                          �   �*  �  �     �     ��. ��<        ������  ����������������        ��d ��                          �   �W  �  �     �     ��. ��=        ������  ����������������        ��d ��  (                        �   0�  �  �     �     ��. ��>        ������  ����������������        ��d ��  2                        �   r�  �  �     �     ��. ��?        ������  ����������������        ��d ��  P                        �    � �  �     �     ��. ��#        ������  ����������������        ��d ��  d                        �   �q �  �     �     ��. ��$        ������  ����������������        ��e ��                          �   �*  �  �     �     ��/ ��@        ������  ����������������        ��e ��                          �   �W  �  �     �     ��/ ��A        ������  ����������������        ��e ��  (                        �   0�  �  �     �     ��/ ��B        ������  ����������������        ��e ��  2                        �   r�  �  �     �     ��/ ��C        ������  ����������������        ��e ��  P                        �    � �  �     �     ��/ ��%        ������  ����������������        ��e ��  d                        �   �q �  �     �     ��/ ��&        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �  �   �� ���        ������  ����������������        ��� ��                            ����    �  �     �     �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �  	  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  
  �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �    �� ���        ������  ����������������        ��� ��                            ����    �  �     �     �� ���        ������  ����������������        ��� ��                            ����    �  �     �  !  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  "  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  #  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  $  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  %  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  &  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  '  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  (  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  )  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  *  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  +  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  ,  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  -  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  .  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  /  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  0  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  1  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  2  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  3  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  4  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  5  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  6  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  7  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  8  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  9  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  :  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  ;  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  <  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  =  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  >  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  ?  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  @  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  A  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  B  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  C  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  D  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  E  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  F  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  G  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  H  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  I  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  J  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  K  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  L  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  M  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  N  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  O  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  P  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  Q  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  R  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  S  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  T  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  U  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  V  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  W  �� ���        ������  ����������������        ��� ��                            ����    �  �     �  X  �� ���        ������  ����������������        ��� ��                            ����    �  �      	  Y  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  Z  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  [  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  \  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  ]  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  ^  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  _  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  `  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  a  �� ���        ������  ����������������        ��� ��                            ����    �  �     		  b  �� ���        ������  ����������������        ��� ��                            ����    �  �     
	  c  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  d  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  e  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  f  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  g  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  h  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  i  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  j  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  k  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  l  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  m  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  n  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  o  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  p  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  q  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  r  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  s  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  t  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  u  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  v  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  w  �� ���        ������  ����������������        ��� ��                            ����    �  �     	  x  �� ���        ������  ����������������        ��� ��                            ����    �  �      	  y  �� ���        ������  ����������������        ��� ��                            ����    �  �     !	  z  �� ���        ������  ����������������        ��� ��                            ����    �  �     "	  {  �� ���        ������  ����������������        ��� ��                            ����    �  �     #	  |  �� ���        ������  ����������������        ��� ��                            ����    �  �     $	  }  �� ���        ������  ����������������        ��� ��                            ����    �  �     %	  ~  �� ���        ������  ����������������        ��� ��                            ����    �  �     &	    �� ���        ������  ����������������        ��� ��                            ����    �  �     '	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     (	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     )	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     *	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     +	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     ,	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     -	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     .	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     /	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     0	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     1	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     2	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     3	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     4	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     5	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     6	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     7	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     8	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     9	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     :	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     ;	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     <	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     =	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     >	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     ?	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     @	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     A	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     B	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     C	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     D	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     E	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     F	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     G	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     H	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     I	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     J	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     K	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     L	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     M	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     N	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     O	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     P	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     Q	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     R	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     S	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     T	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     U	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     V	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     W	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     X	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     Y	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     Z	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     [	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     \	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     ]	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     ^	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     _	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     `	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     a	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     b	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     c	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     d	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     e	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     f	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     g	  �  �� ���        ������  ����������������        ��� ��                            ����    �  �     h	  �  �� ���        ������  ����������������       ����� ��                            �����  �  �    i	      �� ���        ������  ����������������       ����� ��                            �����  �  �    j	      �� ���        ������  ����������������       ����� ��                            �����  �  �    k	      �� ���        ������  ����������������       ����� ��                            �����  �  �    l	      �� ���        ������  ����������������       ����� ��                            �����  �  �    m	      �� ���        ������  ����������������       ����� ��                            �����  �  �    n	      �� ���        ������  ����������������       ����� ��                            �����  �  �    o	      �� ���        ������  ����������������       ����� ��                            �����  �  �    p	      �� ���        ������  ����������������       ����� ��                            �����  �  �    q	      �� ���        ������  ����������������       ����� ��                            �����  �  �    r	      �� ���        ������  ����������������       ����� ��                            �����  �  �    s	      �� ���        ������  ����������������       ����� ��                            �����  �  �    t	      �� ���        ������  ����������������       ����� ��                            �����  �  �    u	      �� ���        ������  ����������������       ����� ��                            �����  �  �    v	      �� ���        ������  ����������������        ��t ��                           ����'   N  �    w	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    x	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    y	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    z	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    {	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    |	      ��X ���        ������  ����������������        ��t ��                           ����'   N  �    }	      ��k ���        ������  ����������������        ��t ��                           ����'   N  �    ~	      ��k ���        ������  ����������������        ��t ��                           ����'   N  �    	      ��l ���        ������  ����������������        ��t ��                           ����'   N  �    �	      ��l ���        ������  ����������������        ��t ��                            ����'   N  �    �	      ��l ���        ������  ����������������        ��d ��  2                        �   '  P�        �	     ��m ���        ������  ����������������        ��e ��  2                        �   '  P�        �	     ��m ���        ������  ����������������       ����� ��                            �����  �        �	     ��l ���        ������  ����������������        ��j ��          h               �����:  `�  �    �	     ��l ���        ������  ����������������       ����� ��                            �����  �        �	     ��l ���        ������  ����������������        ��j ��          h               �����a  �8 �    �	     ��l ���        ������  ����������������        ��i ��                    �     ����    �  �     �	  ~   �� ��>        ������  ����������������        ��i ��                    �     ����    �  �     �	  ~   �� ��>        ������  ����������������        ��i ��        
            �     ����    �  �     �	  ~   �� ��>        ������  ����������������        ��i ��                    �     ����    �  �     �	  ~   �� ��>        ������  ����������������        ��i ���   �             d     ����    �  �     �	     �� ���        ������  ����������������        ��i ���   �             d     ����    �  �     �	     �� ���        ������  ����������������        ��i ���   � 
            d     ����    �  �     �	     �� ���        ������  ����������������        ��i ���   �             d     ����    �  �     �	     �� ���        ������  ����������������        ��i ��   `�              �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   `�              �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   `�  
            �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   `�              �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��                �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��                �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��    
            �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��                �     ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   8 A              �    ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   8 A              �    ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   8 A  
            �    ����    �  �     �	  �   �� ���        ������  ����������������        ��i ��   8 A              �    ����    �  �     �	  �   �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      ��p ���        ������  ����������������       ����� ��                            ����    �  �    �	      ��q ���        ������  ����������������       ����� ��                            ����    �  �    �	      ��r ���        ������  ����������������       ����� ��                            ����    �  �    �	      ��s ���        ������  ����������������       ����� ��                            ����    �  �    �	      ��t ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��T        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��S        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��T        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��S        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��S        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��S        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��V        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��s        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��m        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����   ( 8          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����  ' 5          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����  ' 7          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����  ' 5          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����  ' 7          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������       ����    +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������       ����    +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������       ����    !          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����             � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����             � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����             � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����             � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������       ����    +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����  ! ,          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����   �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������       ����     +          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����    *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����    *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����    *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����    *          � � � d       �  '  P�    �  �	        ���        ������  ����������������       ����    �          2 2 2         �  '  P�    �  �	        ���        ������  ����������������        ��� ��                          ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��                         ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��                         ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��                         ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��                         ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��                          �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��                         �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��                         �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��                         �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��                         �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��                          �����a  P�        �	  �  ��u ���        ������  ����������������        ��� ��   
                      ����P�  ��       �	  �  ��u ���        ������  ����������������        ��� ��                         �����  '        �	  �  ��u ���        ������  ����������������        ��� ��                         �����  '        �	  �  ��u ���        ������  ����������������        ��� ��                         ����'   N        �	      ��u ���        ������  ����������������        ��� ��                        ����'   N        �	      ��u ���        ������  ����������������        ��� ��                        ����'   N        �	      ��u ���        ������  ����������������        ��� ��                        ����'   N        �	      ��u ���        ������  ����������������        ��� ��                        ����'   N        �	      ��u ���        ������  ����������������        ��� ��                         �����:  0u        �	      ��u ���        ������  ����������������        ��� ��                        �����:  0u        �	      ��u ���        ������  ����������������        ��� ��                        �����:  0u        �	      ��u ���        ������  ����������������        ��� ��                        �����:  0u        �	      ��u ���        ������  ����������������        ��� ��                        �����:  0u        �	      ��u ���        ������  ����������������        ��� ��                         �����  '        �	      ��u ���        ������  ����������������        ��� ��                        �����  '        �	      ��u ���        ������  ����������������        ��� ��                        �����  '        �	      ��u ���        ������  ����������������        ��� ��                        �����  '        �	      ��u ���        ������  ����������������        ��� ��   (                      ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��  (                      ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��  (                      ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��  (                      ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��  (                      ����'   N        �	  �  ��u ���        ������  ����������������        ��� ��   F                      �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��  F                      �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��  F                      �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��  F                      �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��  F                      �����:  0u        �	  �  ��u ���        ������  ����������������        ��� ��   Z                      �����  '        �	  �  ��u ���        ������  ����������������        ��� ��  Z                      �����  '        �	  �  ��u ���        ������  ����������������        ��� ��  Z                      �����  '        �	  �  ��u ���        ������  ����������������        ��� ��  Z                      �����  '        �	  �  ��u ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��a        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��b        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��^        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��k        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ���        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��K        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��c        ������  ����������������       ����� ��                            ����    �  �    �	      �� ��d        ������  ����������������       ����� ��                            ����    �  �     
      �� ���        ������
 ����������������       ����� ��                            ����    �  �    
      �� ���        ������ ����������������       ����� ��                            ����    �  �    
      �� ���        ������  ����������������       ����� ��                            ����    �  �    
      �� ��|        ������  ����������������       ����� ��                            ����    �  �    
      �� ��z        ������  ����������������       ����� ��                            ����    �  �    
      �� ���        ������  ����������������       ����� ��                            ����    �  �    
      �� ��q        ������  ����������������       ����� ��                            ����    �  �    
      �� ���        ������  ����������������       ����� ��                            ����    �  �    
      �� ���        ������  ����������������       ����� ��                            ����    �  �    	
      �� ���        ������  ����������������       ����� ��                            ����    �  �    

      �� ��l        ������  ����������������       ����� ��                            ����    �  �    
      �� ��        ������  ����������������       ����� ��                            ����    �  �    
      �� ���        ������  ����������������        ��� ��                           ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                          ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                          ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                          ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                          ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                          ����    �  �     
  �   �� ���        ������  ����������������        ��� ��                         ����    �  �     
  �   �� ���        ������  ����������������        ��� ��#                       ����    �  �     
  �   �� ���        ������  ����������������        ��� ��# (                      ����    �  �     
  �   �� ���        ������  ����������������        ��� ��$                       ����    �  �     
  �   �� ���        ������  ����������������        ��� ��$ (                      ����    �  �     
  �   �� ���        ������  ����������������        ��t ��            #               ������ ���      
      �� ��	        ������  ����������������        ��� ��)                       ����    �  �     s
  �   �� ���        ������  ����������������        ��� ��)                       ����    �  �     t
  �   �� ���        ������  ����������������        ��� ��)     
                  ����    �  �     u
  �   �� ���        ������  ����������������        ��� ��& d   <                    ����    �  �     v
  h   �� ���        ������  ����������������        ��� ��& d   <  
                  ����    �  �     w
  h   �� ���        ������  ����������������        ��� ��& d   <                    ����    �  �     x
  h   �� ���        ������  ����������������        ��� ��& d   <                    ����    �  �     y
  h   �� ���        ������  ����������������        ��� ��& d   x                    ����    �  �     z
  h   �� ���        ������  ����������������        ��� ��& d   x  
                  ����    �  �     {
  h   �� ���        ������  ����������������        ��� ��& d   x                    ����    �  �     |
  h   �� ���        ������  ����������������        ��� ��& d   x                    ����    �  �     }
  h   �� ���        ������  ����������������        ��d ��  P                        �       �  �     ~
     ��. ��#        ������  ����������������        ��d ��  d                        �       �  �     
     ��. ��$        ������  ����������������        ��e ��  P                        �       �  �     �
     ��/ ��%        ������  ����������������        ��e ��  d                        �       �  �     �
     ��/ ��&        ������  ����������������        ���  -     ,                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  -     X                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  -     �                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  -     `	                   ����    �  �     �
  �   �� ���        ������  ����������������       ����� ��                            ������� `*�     �
      �� ���        ������  ����������������       ����� ��                            ���� ����#    �
      �� ���        ������  ����������������        ���  .     ,                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  .     X                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  .     �                   ����    �  �     �
  �   �� ���        ������  ����������������        ���  .     `	                   ����    �  �     �
  �   �� ���        ������  ����������������        ��� ��                           ����    �  �     �
  �   �� ���        ������  ����������������        ��� ��         
                  ����    �  �     �
  �   �� ���        ������  ����������������        ��� ��                           ����    �  �     �
  �   �� ���        ������  ����������������        ��� ��                           ����    �  �     �
  �   �� ���        ������  ����������������        ��i ���   �                   ����    '  �     �
  �   �� ��>        ������  ����������������        ��i ���   �                   ����    '  �     �
  �   �� ��>        ������  ����������������        ��i ���   �                   ����    '  �     �
  �   �� ��>        ������  ����������������        ��t ��            $               ����'   N       �
      �� ��R        ������  ����������������          ����	y
�2    Io���     ~4  v 8�   ��  �
      �    �    ������� � �����  �  �            ����	�
�2    Rw���     �4  � ��   ��  �
     �    �    ������� � �����  �  �            ����	�
�2    [���     b5  �
 H�   ��  �
     �    �    ������� � �����  �  �            ��	 
�
2    d����     �5  $ �   ��  �
     �    �   ������� � �����  �  �            ��)	G
$B2    m����     F6  ^ X3   ��  �
     �    �   ������� �����  �  �            ��O	n
On2    v����     �6  � �_   ��  �
     �    �   ������� �����  �  �            ��u	�
z�2    ����     *7  � h�   ��  �
     �    �   ������� �����  �  �            ���	�
��2    �����     �7   �   ��  �
     �    �   ������� �����  �  �            ���	�
��2    �����     8  F x�   ��  �
     �    �   ������� �����  �  �            ���	
�2    �����     �8  �     ��  �
	     �    �   ������� &)   �  �  �            ��%��
2    Io���     2=  h# ��   ��  �
      �    �    ������� � �����  �  �            ��V��C2    Rw���     �=  �% �   ��  �
     �    �    ������� � �����  �  �            ����}2    [���     .>  ( �I   ��  �
     �    �    ������� � �����  �  �            ���*D�2    d����     �>  p* 0{   ��  �
     �    �   ������� � �����  �  �            ���]|�2    m����     *?  �, h�   ��  �
     �    �   ������� �����  �  �            ����)2    v����     �?   / ��   ��  �
     �    �   ������� �����  �  �            ��K��c2    ����     &@  x1 �   ��  �
     �    �   ������� �����  �  �            ��|�#�2    �����     �@  �3 @   ��  �
     �    �   ������� �����  �  �            ���'[�2    �����     "A  (6 Hq   ��  �
     �    �   ������� �����  �  �            ���Z�2    �����     �A  �8 ��   ��  �
	     �    �   ������� &�����  �  �            �����2    X~���     �4  f ��   ��  �
      �   �    ������� � �����  �  �            ������2    a����      5  �	 ��   ��  �
     �   �    ������� � �����  �  �            �����	2    j����     �5  � �   ��  �
     �   �    ������� � �����  �  �            ��,	2    s����     6   �   ��  �
     �   �   ������� � �����  �  �            ��5F%P	2    |����     v6  N F   ��  �
     �   �   ������� �����  �  �            ��cuHu	2    �����     �6  � �r   ��  �
     �   �   ������� �����  �  �            ����k�	2    �����     Z7  � (�   ��  �
     �   �   ������� �����  �  �            ������	2    �����     �7  � ��   ��  �
     �   �   ������� �����  �  �            �����	2    �����     >8  6 8�   ��  �
     �   �   ������� �����  �  �            ��0�
2    �����     �8  p �$   ��  �
	     �   �   ������� &[   �  �  �            ���N�	^2    X~���     d=  X$ 8�   ��  �
      �   �    ������� � �����  �  �            ��-�
�2    a����     �=  �& p,   ��  �
     �   �    ������� � �����  �  �            ��h�<
�2    j����     `>  ) �]   ��  �
     �   �    ������� � �����  �  �            ���i
�2    s����     �>  `+ ��   ��  �
     �   �   ������� � �����  �  �            ���B�
2    |����     \?  �- �   ��  �
     �   �   ������� �����  �  �            ���
K2    �����     �?  0 P�   ��  �
     �   �   ������� �����  �  �            ��U��
z2    �����     X@  h2 �"   ��  �
     �   �   ������� �����  �  �            ���� �2    �����     �@  �4 �S   ��  �
     �   �   ������� �����  �  �            ���5M�2    �����     TA  7 ��   ��  �
     �   �   ������� �����  �  �            ��r{2    �����     �A  p9 0�   ��  �
	     �   �   ������� &�����  �  �            ���	�
�	�
2    �����     �4  � �   ��  �
      �   �    ������� � �����  �  �            ���	�
�	�
2    ���     �4  � p�   ��  �
     �   �    ������� � �����  �  �            ���	�	2    ���     n5  & ��   ��  �
     �   �    ������� � �����  �  �            ��
/
/2    ���     �5  ` �   ��  �
     �   �   ������� � �����  �  �            ��:
X:
X2    #�#��     R6  � 8   ��  �
     �   �   ������� �����  �  �            ��c
�c
�2    ,�,��     �6  � �d   ��  �
     �   �   ������� �����  �  �            ���
��
�2    5�5��     67   �   ��  �
     �   �   ������� �����  �  �            ���
��
�2    >�>��     �7  H ��   ��  �
     �   �   ������� �����  �  �            ���
��
�2    G�G��     8  � (�   ��  �
     �   �   ������� �����  �  �            ��((2    PP��     �8  � �   ��  �
	     �   �   ������� &�   �  �  �            ��z�z�2    �����     >=  �# t�   ��  �
      �   �    ������� � �����  �  �            ����2    ���     �=  �% �   ��  �
     �   �    ������� � �����  �  �            ���S�S2    ���     :>  T( �N   ��  �
     �   �    ������� � �����  �  �            ����2    ���     �>  �* �   ��  �
     �   �   ������� � �����  �  �            ��L�L�2    #�#��     6?  - T�   ��  �
     �   �   ������� �����  �  �            ������2    ,�,��     �?  \/ ��   ��  �
     �   �   ������� �����  �  �            ���,�,2    5�5��     2@  �1 �   ��  �
     �   �   ������� �����  �  �            ���b�b2    >�>��     �@  4 �D   ��  �
     �   �   ������� �����  �  �            ����2    G�G��     .A  d6 4v   ��  �
     �   �   ������� �����  �  �            ��R�R�2    PP��     �A  �8 l�   ��  �
	     �   �   ������� &�����  �  �            ��y
���	2    Sy���     �4  * H�   ��  �
      �   �    ������� � �����  �  �            ���
���	2    \����     5  d	 л   ��  �
     �   �    ������� � �����  �  �            ���
���	2    e����     �5  � X�   ��  �
     �   �    ������� � �����  �  �            ���
	 
2    n����     �5  � �   ��  �
     �   �   ������� � �����  �  �            ��$B)	G
2    w����     j6   hA   ��  �
     �   �   ������� �����  �  �            ��OnO	n
2    �����     �6  L �m   ��  �
     �   �   ������� �����  �  �            ��z�u	�
2    �����     N7  � x�   ��  �
     �   �   ������� �����  �  �            �����	�
2    �����     �7  �  �   ��  �
     �   �   ������� �����  �  �            �����	�
2    �����     28  � ��   ��  �
     �   �   ������� �����  �  �            ����	
2    �����     �8  4     ��  �
	     �   �   ������� &�   �  �  �            ���
%�2    Sy���     W=  $ L�   ��  �
         �    ������� � �����  �  �            ���CV�2    \����     �=  t& �'   ��  �
        �    ������� � �����  �  �            ��}��2    e����     S>  �( �X   ��  �
        �    ������� � �����  �  �            ��D��*2    n����     �>  $+ �   ��  �
        �   ������� � �����  �  �            ��|��]2    w����     O?  |- ,�   ��  �
        �   ������� �����  �  �            ���)�2    �����     �?  �/ d�   ��  �
        �   ������� �����  �  �            ���cK�2    �����     K@  ,2 �   ��  �
        �   ������� �����  �  �            ��#�|�2    �����     �@  �4 �N   ��  �
        �   ������� �����  �  �            ��[��'2    �����     GA  �6 �   ��  �
        �   ������� �����  �  �            ����Z2    �����     �A  49 D�   ��  �
	        �   ������� &�����  �  �            �����2    �QN��     r4  : �|   ��  �
        �    ������� � �����  �  �            ������2    �YW��     �4  t �   ��  �
       �    ������� � �����  �  �            ���	��2    �a`��     V5  �
 ��   ��  �
       �    ������� � �����  �  �            ��,	2    �ii��     �5  �     ��  �
       �   ������� � �����  �  �            ��%P	5F2    �qr��     :6  " �.   ��  �
       �   ������� �����  �  �            ��Hu	cu2    y{��     �6  \ 0[   ��  �
       �   ������� �����  �  �            ��k�	��2    ����     7  � ��   ��  �
       �   ������� �����  �  �            ����	��2    ����     �7  � @�   ��  �
       �   ������� �����  �  �            ����	�2    ����     8  
 ��   ��  �
       �   ������� �����  �  �            ���
02    "����     t8  D P   ��  �
	       �   ������� &�   �  �  �            ���	^�N2    �QN��     %=  ,# ��   ��  �
        �    ������� � �����  �  �            ��
�-�2    �YW��     �=  �% �   ��  �
       �    ������� � �����  �  �            ��<
�h�2    �a`��     !>  �' E   ��  �
       �    ������� � �����  �  �            ��i
��2    �ii��     �>  4* Dv   ��  �
       �   ������� � �����  �  �            ���
�B2    �qr��     ?  �, |�   ��  �
       �   ������� �����  �  �            ���
K2    y{��     �?  �. ��   ��  �
       �   ������� �����  �  �            ���
zU�2    ����     @  <1 �	   ��  �
       �   ������� �����  �  �            �� ���2    ����     �@  �3 $;   ��  �
       �   ������� �����  �  �            ��M��52    ����     A  �5 \l   ��  �
       �   ������� �����  �  �            ��{r2    "����     �A  D8 ��   ��  �
	       �   ������� &�����  �  �             		"
		"

2    �����     �4  � ��   ��  �
        �    ������� � �����  �  �             0	J
0	J

2    ���     5  (	  �   ��  �
       �    ������� � �����  �  �             W	r
W	r

2    ���     z5  b ��   ��  �
       �    ������� � �����  �  �             ~	�
~	�

2    ���     �5  � 0   ��  �
       �   ������� � �����  �  �             �	�
�	�

2    !�#��     ^6  � �<   ��  �
       �   ������� �����  �  �             �	�
�	�

2    *�,��     �6   @i   ��  �
       �   ������� �����  �  �             �	�	
2    3�5��     B7  J ȕ   ��  �
       �   ������� �����  �  �             
<
<
2    <�>��     �7  � P�   ��  �
       �   ������� �����  �  �             A
dA
d
2    E�G��     &8  � ��   ��  �
       �   ������� �����  �  �             h
�h
�
2    NP��     �8  � `   ��  �
	       �   ������� &#  �  �  �             �,�,
2    �����     K=  �# `�   ��  �
        �    ������� � �����  �  �             �`�`
2    ���     �=  8& �"   ��  �
       �    ������� � �����  �  �             $�$�
2    ���     G>  �( �S   ��  �
       �    ������� � �����  �  �             W�W�
2    ���     �>  �* �   ��  �
       �   ������� � �����  �  �             ����
2    !�#��     C?  @- @�   ��  �
       �   ������� �����  �  �             �2�2
2    *�,��     �?  �/ x�   ��  �
       �   ������� �����  �  �             �f�f
2    3�5��     ?@  �1 �   ��  �
       �   ������� �����  �  �             !�!�
2    <�>��     �@  H4 �I   ��  �
       �   ������� �����  �  �             T�T�
2    E�G��     ;A  �6  {   ��  �
       �   ������� �����  �  �             ��
2    NP��     �A  �8 X�   ��  �
	       �   ������� &�����  �  �             �
��2    �%���     �4  f ��   ��  �
        �    ������� � �����  �  �             G��2    �.���      5  �	 ��   ��  �
       �    ������� � �����  �  �             @u�	2    �7���     �5  � �   ��  �
       �    ������� � �����  �  �             l�,	2    �@���     6   �   ��  �
       �   ������� � �����  �  �             ��%P	2    �I���     v6  N F   ��  �
       �   ������� �����  �  �             ��Hu	2    �R���     �6  � �r   ��  �
       �   ������� �����  �  �             �+k�	2    �[���     Z7  � (�   ��  �
       �   ������� �����  �  �             X��	2    �d���     �7  � ��   ��  �
       �   ������� �����  �  �             I���	2    �m���     >8  6 8�   ��  �
       �   ������� �����  �  �             u��
2    �v���     �8  p �$   ��  �
	       �   ������� &)   �  �  �             ����2    �%���     d=  X$ 8�   ��  �
        �    ������� � �����  �  �             f�
�2    �.���     �=  �& p,   ��  �
       �    ������� � �����  �  �             �2<
�2    �7���     `>  ) �]   ��  �
       �    ������� � �����  �  �             �mi
�2    �@���     �>  `+ ��   ��  �
       �   ������� � �����  �  �             ��
2    �I���     \?  �- �   ��  �
       �   ������� �����  �  �             L��
K2    �R���     �?  0 P�   ��  �
       �   ������� �����  �  �             ��
z2    �[���     X@  h2 �"   ��  �
       �   ������� �����  �  �             �Y �2    �d���     �@  �4 �S   ��  �
       �   ������� �����  �  �             ��M�2    �m���     TA  7 ��   ��  �
       �   ������� �����  �  �             2�{2    �v���     �A  p9 0�   ��  �
	       �   ������� &�����  �  �           ��q  � � � �  �    � � D v d     �   t  �1        �
      �� ���        ������  ����������������         ��q  KQKQ �    Q � �     �   8  ��        �
      �� ���        ������  ����������������        ��� �� d                       �     �     �
  �  �� ���        ������  ����������������        ��� �� d                       �     �     �
  �  �� ���        ������  ����������������        ��� �� d                       �     �     �
     �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d                       �     �     �
  	  �� ���        ������  ����������������        ��� �� d  m                    �     �     �
  
  �� ���        ������  ����������������        ��� �� d                       �     �     �
    �� ���        ������  ����������������        ��� �� d   
                     �     �     �
    �� ���        ������  ����������������        ��� ��                        ��     �     �
    �� ���        ������  ����������������        ��� ��                         ��     �     �
    �� ���        ������  ����������������        ��� ��                     ��     �     �
    �� ���        ������  ����������������        ��� ��                       ��     �     �
    �� ���        ������  ����������������        ��� ��     
                 ��     �     �
    �� ���        ������  ����������������        ��� �� 
 
                     �      �     �
    �� ���        ������  ����������������        ��� �� 
 
                     �      �     �
    �� ���        ������  ����������������        ��� �� 
 
   
                  '      �     �
    �� ���        ������  ����������������        ��� ��                        ��     �     �
    �� ���        ������  ����������������        ��� ��                          ��     �     �
    �� ���        ������  ����������������        ��� ��                           ����'  P�        �
    ��9 ���        ������ ����������������        ��� ��                           ���� N  P�        �
    ��9 ���        ������( ����������������        ��� ��                           ����@�  P�        �
    ��9 ���        ������< ����������������        ��� ��                           �����8 P�        �
    ��9 ���        ������P ����������������        ��� ��                           ���� q P�        �
    ��9 ���        ������x ����������������        ��� ��                           ���� q P�        �
    ��9 ���        ������� ����������������        ��� ��                           ����'  P�        �
    ��x ���        ������ ����������������        ��� ��                           ���� N  P�        �
    ��x ���        ������* ����������������        ��� ��                           ����@�  P�        �
    ��x ���        ������6 ����������������        ��� ��                           �����8 P�        �
    ��x ���        ������K ����������������        ��� ��                           ���� q P�        �
    ��x ���        ������� ����������������        ��� ��                           ���� q P�        �
    ��x ���        ������� ����������������        ���                              ����'  P�        �
    ��x ���        ������ ����������������        ��� *                             ����'  P�        �
    ��x ���        ������ ����������������        ���                              ����0u  P�        �
    ��x ���        ������P ����������������        ���                              ����0u  P�        �
    ��x ���        ������P ����������������        ��� 0                             ����0u  P�        �
    ��x ���        ������P ����������������        ���                              ����P�  P�        �
    ��x ���        ������n ����������������        ���                              ����P�  P�        �
    ��x ���        ������n ����������������        ���                              ����P�  P�        �
    ��x ���        ������n ����������������        ���                              ����P�  P�        �
    ��x ���        ������n ����������������        ���                              ����P�  P�        �
    ��x ���        ������n ����������������        ���                               ����P�  P�        �
    ��x ���        ������n ����������������        ��� ��         
                  ����'  �� �     �
    �� ���        ������������������������        ��� ��                           ����PF   � �     �
    �� ���        ������������������������        ��� ��                           �����a  �� �     �
    �� ���        ������������������������        ��� ��                            �����  �  �     �
    �� ���        ������������������������        ��� ��                            �����  �  �     �
    �� ���        ������������������������        ��� ��                            ����@  @  �     �
    �� ���        ������������������������          ��*�"2    �6� �       '  �t  P�        
         �     �m�    �    �  �  �             ��c�l2    �<� �       U  �u  ��                 �     �m�    �    �  �  �             ���X�2    �B� �       �  `w  �                 �     �m�    �    �  �  �             ���]�(2    �H� �       �  �x  ("                 �     �m�    �    �  �  �             ��:��2    �N� �       �  0z  p4                 �     �m�    �    �  �  �             ����l�2    �T� �         �{  �F                 �     �m�    �    �  �  �             ���U�2    �S� �         �  8p        
         �    TX�       �  �  �             ���M�2    �Y� �       A  ��  ��                 �    TX�       �  �  �             ��*��i2    �_� �       x  �  ��                 �    TX�       �  �  �             ���h�2    e� �       �  ��  4�                 �    TX�       �  �  �             ���]�O2    k� �       �  �  ��                 �    TX�       �  �  �             ��3�1�2    q� �         ��  ��                 �    TX�       �  �  �             ����]2    z� �       �  ��  �2	   ��   
         �    :��    �    �  �  �             ��f�E�2    "�� �       �  ��  ~K	   ��            �    :��    �    �  �  �             ���7�$2    *�� �       
  F�  d	   ��            �    :��    �    �  �  �             ��!�%�2    2�� �       I  �  �|	   ��            �    :��    �    �  �  �             ��}�*2    :��       �  ��  R�	   ��            �    :��    �    �  �  �             ����	�2    B��       �  2�  �	   ��            �    :��    �    �  �  �             ���&�2    H�      �  ~�  �7   ��   
         �    �Z       �  �  �             ������2    P�         @�   T   ��            �    �Z       �  �  �             ��U�b�2    X�      H  �   p   ��            �    �Z       �  �  �             ���l��2    `�       �  ĸ  @�   ��            �    �Z       �  �  �             ��9�r!2    h�&      �  ��  `�   ��            �    �Z    
   �  �  �             ���[��2    p�,          H�  ��   ��            �    �Z    	   �  �  �             ��4�=�2    u�."n     �"  ��  ă   ��   
         �   ���       �  �  �            ���&�F2    }�4(o     �"  d�  ��   ��            �   ���       �  �  �            ����%�2    ��:.p     <#  D�  ��   ��            �   ���       �  �  �            ��~+�|2    ��@4q     �#  $�  d�   ��            �   ���       �  �  �            ����U	2    ��F:r     �#  �  D   ��            �   ���       �  �  �            ��o5��	2    ��L@s     0$  ��  $#   ��            �   ���       �  �  �            ���h��2    ��MAx     ;)  �      ��   
         �   ���       �  �  �            ��,�t2    ��SGy     �)  �  �>   ��            �   ���       �  �  �            ���V��2    ��YMz     �)  �  �b   ��            �   ���       �  �  �            ��2��r	2    ��_S{     N*  
�  ��   ��            �   ���       �  �  �            ����M	
2    �eY|     �*  �  ��   ��            �   ���       �  �  �            ��='	�	�
2    �k_}     +  �  l�   ��            �   ���       �  �  �            ��d�k2    �l`�     �0  "  �   ��   
            ���    	    �  �  �            ����>	2    �rf�     1  > �*   ��               ���    !   �  �  �            ��Q"��	2    �'xl�     w1  Z �R   ��               ���    "   �  �  �            �����	�
2    �/~r�     �1  v �z   ��               ���    #   �  �  �            ���|	J
=2    7�x�     D2  � ֢   ��               ���    $   �  �  �            ��"	&
2    ?�~�     �2  �
 ��   ��               ���    %   �  �  �            ��	��C	2    D���     �8  � �>   ��   
         '   ���    $    �  �  �            ���a	�	2    L���     d9  � k   ��            '   ���    /!   �  �  �            ����	�
2    &T���     �9  .! ��   ��            '   ���    ."   �  �  �            ����	�
�2    /\���     H:  h#  �   ��            '   ���    -#   �  �  �            ��e	t
[^2    8d���     �:  �% ��   ��            '   ���    ,$   �  �  �            ��
0&<2    Al���     ,;  �' 0   ��            '   ���    +%   �  �  �            ����W	'
2    Gp���     B  �: ��   ��   
         (   ���    *   �  �  �            ��C.	�	�
2    Px���     �B  0= �   ��            (   ���    +   �  �  �            ����	�
�2    Y����     C  �? (6   ��            (   ���    
,   �  �  �            ���	�
��2    b����     �C  �A `g   ��            (   ���    	-   �  �  �            ��O
ux�2    k����     D  8D ��   ��            (   ���    .   �  �  �            ��BX�2    t����     �D  �F ��   ��            (   ���    /   �  �  �            ��)
ASX2    ����     �8  � �>   ��  �

     �    �   ���    %*   �  �  �            ���
/G2    ����     d9  � k   ��  �
     �    �   ���    $+   �  �  �            ����G2    ���     �9  .! ��   ��  �
     �    �   ���    #,   �  �  �            ���a�2    ���     H:  h#  �   ��  �
     �    �   ���    "-   �  �  �            ���t�2    �� �     �:  �% ��   ��  �
     �    �   ���    !.   �  �  �            ����2    ��'�     ,;  �' 0   ��  �
     �    �   ���     /   �  �  �            ��Q���2    ����     B  �: ��   ��  �

     �    �   ���    %*   �  �  �            ��z��2    ����     �B  0= �   ��  �
     �    �   ���    $+   �  �  �            ���l�2    ���     C  �? (6   ��  �
     �    �   ���    #,   �  �  �            �� �-�2    ���     �C  �A `g   ��  �
     �    �   ���    "-   �  �  �            ���a�2    �� �     D  8D ��   ��  �
     �    �   ���    !.   �  �  �            ��+��I2    ��'�     �D  �F ��   ��  �
     �    �   ���     /   �  �  �            ��r�82    �E� �       F  �u  ��       # 
     !   �    �}Y    � 4   �  �  �             ��[�r2    �K� �       u  �v  �	       #      !   �    �}Y    � 5   �  �  �             ���C�2    �Q� �       �  Px         #      !   �    �}Y    � 6   �  �  �             ����2    �W� �       �  �y  X.       #      !   �    �}Y    � 7   �  �  �             ��p��M2    �]� �          {  �@       #      !   �    �}Y    � 8   �  �  �             ���[�2    �c� �       1  �|  �R       #      !   �    �}Y    � 9   �  �  �             ���I�2    �b� �       +  �  X}       $ 
     "   �    P�b    4   �  �  �             ��x��2    h� �       a  z�  ��       $      "   �    P�b    5   �  �  �             ��\��A2    
n� �       �   �   �       $      "   �    P�b    6   �  �  �             ���`�2    t� �       �  ��  T�       $      "   �    P�b    7   �  �  �             ��@�c�2    z� �         �  ��       $      "   �    P�b    8   �  �  �             ���M�N2    "�� �       9  ��  ��       $      "   �    P�b    9   �  �  �             ��N��42    )�� �       �  �  �@	   ��  % 
     #   �    66�    � >   �  �  �             ���4�2    1�� �       �  ��  �Y	   ��  %      #   �    66�    � ?   �  �  �             ���B�2    9�� �       .  6�  *r	   ��  %      #   �    66�    � @   �  �  �             ���=�?2    A�� �       m  ڢ  Ɗ	   ��  %      #   �    66�    � A   �  �  �             �����2    I��       �  ~�  b�	   ��  %      #   �    66�    � B   �  �  �             ���IP2    Q��       �  "�  ��	   ��  %      #   �    66�    � C   �  �  �             ���0�2    W�      �  n�  �F   ��  & 
     $   �    ��    >   �  �  �             ��m {2    _�      &  0�   c   ��  &      $   �    ��    ?   �  �  �             ���~�i2    g�      n  �      ��  &      $   �    ��    @   �  �  �             ��*9�2    o�       �  ��  @�   ��  &      $   �    ��    A   �  �  �             ����O2    w�&      �  v�  `�   ��  &      $   �    ��    
B   �  �  �             ���Y	��2    �,       F  8�  ��   ��  &      $   �    ��    	C   �  �  �             ���V�J2    ��."n     �"  t�  ��   ��  ' 
     %   �   ���    H   �  �  �            ��7���2    ��4(o     #  T�  ��   ��  '      %   �   ���    I   �  �  �            ���fW2    ��:.p     f#  4�  t�   ��  '      %   �   ���    J   �  �  �            ��j'	��2    ��@4q     �#  �  T�   ��  '      %   �   ���    K   �  �  �            ��	�	:2    ��F:r     
$  ��  4   ��  '      %   �   ���    L   �  �  �            ���	{
��2    ��L@s     \$  ��  3   ��  '      %   �   ���    M   �  �  �            ���2/�2    ��MAx     f)   �   ,   ��  ( 
     &   �   ���    H   �  �  �            ����H2    ��SGy     �)  ��  �O   ��  (      &   �   ���    I   �  �  �            ���a	��2    �YMz     *  ��  �s   ��  (      &   �   ���    J   �  �  �            ��i	:
yS2    �_S{     z*  ��  ��   ��  (      &   �   ���    K   �  �  �            ��
�
��2    �eY|     �*  ��  p�   ��  (      &   �   ���    L   �  �  �            ���
�ic2    �k_}     2+  ��  L�   ��  (      &   �   ���    M   �  �  �            ��^	�z2    �&l`�     �0   V   ��  ) 
     '      ���    	R   �  �  �            ����	$�2    �.rf�     ?1  . j<   ��  )      '      ���    S   �  �  �            ���	m
�k2    6xl�     �1  J ~d   ��  )      '      ���    T   �  �  �            ��q
]*2    
>~r�     2  f ��   ��  )      '      ���    U   �  �  �            ��,)��2    F�x�     t2  �	 ��   ��  )      '      ���    V   �  �  �            ���3A	2    N�~�     �2  � ��   ��  )      '      ���    W   �  �  �            ��>		
N$2    #S���     "9  � HQ   ��  * 
     (   )   ���    $R   �  �  �            ���	�
��2    ,[���     �9  � �}   ��  *      (   )   ���    /S   �  �  �            ���
}8-2    5c���     :  " X�   ��  *      (   )   ���    .T   �  �  �            ������2    >k���     x:  X$ ��   ��  *      (   )   ���    -U   �  �  �            ��Wfk�	2    Gs���     �:  �& h   ��  *      (   )   ���    ,V   �  �  �            ��4V	4
2    P{���     \;  �( �/   ��  *      (   )   ���    +W   �  �  �            ��'
��2    V���     PB  �; h�   ��  + 
     )   *   ���    \   �  �  �            ���
�g[2    _����     �B   > �   ��  +      )   *   ���    ]   �  �  �            ������2    h����     LC  x@ �I   ��  +      )   *   ���    
^   �  �  �            ������	2    q����     �C  �B {   ��  +      )   *   ���    	_   �  �  �            ����=	m
2    z����     HD  (E H�   ��  +      )   *   ���    `   �  �  �            �����	(2    �����     �D  �G ��   ��  +      )   *   ���    a   �  �  �            ��hy	5
2    ����     "9  � HQ   ��  �

     �   �   ���    %\   �  �  �            ��X|�	�
2    ����     �9  � �}   ��  �
     �   �   ���    $]   �  �  �            ��Y�f
�2    ���     :  " X�   ��  �
     �   �   ���    #^   �  �  �            ���V�2    ���     x:  X$ ��   ��  �
     �   �   ���    "_   �  �  �            ���S!�2    �� �     �:  �& h   ��  �
     �   �   ���    !`   �  �  �            ��(���2    ��'�     \;  �( �/   ��  �
     �   �   ���     a   �  �  �            ��n�	9
2    ����     PB  �; h�   ��  �

     �   �   ���    %\   �  �  �            ��^��	�
2    ����     �B   > �   ��  �
     �   �   ���    $]   �  �  �            ��`�k
�2    ���     LC  x@ �I   ��  �
     �   �   ���    #^   �  �  �            ���[�2    ���     �C  �B {   ��  �
     �   �   ���    "_   �  �  �            ���]'�2    �� �     HD  (E H�   ��  �
     �   �   ���    !`   �  �  �            ��0� �2    ��'�     �D  �G ��   ��  �
     �   �   ���     a   �  �  �            ��{�{�2    �� ��       /  �t  \�       7 
     5   �    �V#    � f   �  �  �             ��� � 2    �� ��       ^  4v  �        7      5   �    �V#    � g   �  �  �             ���j�j2    �� ��       �  �w  �       7      5   �    �V#    � h   �  �  �             ��X�X�2    �� ��       �  y  4%       7      5   �    �V#    � i   �  �  �             ���&�&2    �� ��       �  lz  |7       7      5   �    �V#    � j   �  �  �             ������2    �� ��         �{  �I       7      5   �    �V#    � k   �  �  �             ���i�i2    �� ��         @�  �s       8 
     6   �    ��H    f   �  �  �             ��B�B�2    �� ��       H  Ɖ  Ԉ       8      6   �    ��H    g   �  �  �             ����2    �� ��       ~  L�  (�       8      6   �    ��H    h   �  �  �             ������2    �� ��       �  Ҍ  |�       8      6   �    ��H    i   �  �  �             ��P�P�2    �� ��       �  X�  ��       8      6   �    ��H    j   �  �  �             ���M�M2    �� ��          ޏ  $�       8      6   �    ��H    k   �  �  �             ����2    �� ��       �  :�  f6	   ��  9 
     7   �    <|�    � p   �  �  �             ���`�`2    �� ��       �  ޞ  O	   ��  9      7   �    <|�    � q   �  �  �             ��1�1�2    � ��         ��  �g	   ��  9      7   �    <|�    � r   �  �  �             ���E�E2    ���       R  &�  :�	   ��  9      7   �    <|�    � s   �  �  �             ����2    �
��       �  ʣ  ֘	   ��  9      7   �    <|�    � t   �  �  �             ��z-z-2    ��      �  n�  r�	   ��  9      7   �    <|�    � u   �  �  �             ����2    
      �  ��  �;   ��  : 
     8   �    ׂ�    p   �  �  �             ��yy2          	  |�  �W   ��  :      8   �    ׂ�    q   �  �  �             ���y�y2    "      Q  >�  �s   ��  :      8   �    ׂ�    r   �  �  �             ��bb2     (       �   �   �   ��  :      8   �    ׂ�    s   �  �  �             ������2    (.("      �  º   �   ��  :      8   �    ׂ�    
t   �  �  �             ��OO2    040(      )  ��  @�   ��  :      8   �    ׂ�    	u   �  �  �             ���X�X2    666*n     �"  ��  ��   ��  ; 
     9   �   ���    z   �  �  �            ��&�&�2    ><>0o     �"  ��  ��   ��  ;      9   �   ���    {   �  �  �            ���C�C2    FBF6p     D#  ��  ��   ��  ;      9   �   ���    |   �  �  �            ��+�+�2    NHN<q     �#  `�  `�   ��  ;      9   �   ���    }   �  �  �            ���x�x2    VNVBr     �#  @�  @   ��  ;      9   �   ���    ~   �  �  �            ��5	5	2    ^T^Hs     7$   �   '   ��  ;      9   �   ���       �  �  �            ��dd2    cUcIx     F)  L�  X   ��  < 
     :   �   ���    z   �  �  �            ������2    k[kOy     �)  J�  4C   ��  <      :   �   ���    {   �  �  �            ��QQ2    sasUz     �)  H�  g   ��  <      :   �   ���    |   �  �  �            ������2    {g{[{     Z*  F�  �   ��  <      :   �   ���    }   �  �  �            ���d	�d	2    �m�a|     �*  D�  Ȯ   ��  <      :   �   ���    ~   �  �  �            ��"	
"	
2    �s�g}     +  B�  ��   ��  <      :   �   ���       �  �  �            ����2    �t�h�     �0  ^  �   ��  = 
     ;      ���    	�   �  �  �            ���V�V2    �z�n�     1  z /   ��  =      ;      ���    �   �  �  �            ����2    ���t�     �1  � "W   ��  =      ;      ���    �   �  �  �            ����	��	2    ���z�     �1  � 6   ��  =      ;      ���    �   �  �  �            ��v	g
v	g
2    �����     R2  � J�   ��  =      ;      ���    �   �  �  �            �� 
" 
"2    �����     �2  �
 ^�   ��  =      ;      ���    �   �  �  �            ������2    �����     �8  � 8C   ��  > 
     <   +   ���    $�   �  �  �            ��[5	[5	2    �����     p9  0 �o   ��  >      <   +   ���    /�   �  �  �            ����	��	2    �����     �9  j! H�   ��  >      <   +   ���    .�   �  �  �            ���	�
�	�
2    �����     T:  �# ��   ��  >      <   +   ���    -�   �  �  �            ��m
~m
~2    �����     �:  �% X�   ��  >      <   +   ���    ,�   �  �  �            ��(L(L2    �����     8;  ( �!   ��  >      <   +   ���    +�   �  �  �            ���m	�m	2    �����     *B  ; ��   ��  ? 
     =   ,   ���    �   �  �  �            ��,	
,	
2    ���     �B  l= �	   ��  ?      =   ,   ���    �   �  �  �            ���	�
�	�
2    ���     &C  �? ;   ��  ?      =   ,   ���    
�   �  �  �            ���
��
�2    ���     �C  B Ll   ��  ?      =   ,   ���    	�   �  �  �            ��s�s�2    ���     "D  tD ��   ��  ?      =   ,   ���    �   �  �  �            ��@x@x2    '�'��     �D  �F ��   ��  ?      =   ,   ���    �   �  �  �            ��I^I^2    YY �     �8  � 8C   ��  �

     �   �   ���    %�   �  �  �            ��<<2    bb�     p9  0 �o   ��  �
     �   �   ���    $�   �  �  �            ���)�)2    kk�     �9  j! H�   ��  �
     �   �   ���    #�   �  �  �            ��oo2    t!t�     T:  �# ��   ��  �
     �   �   ���    "�   �  �  �            ����2    }(}�     �:  �% X�   ��  �
     �   �   ���    !�   �  �  �            ����2    �/�#�     8;  ( �!   ��  �
     �   �   ���     �   �  �  �            ��NbNb2    YY �     *B  ; ��   ��  �

     �   �   ���    %�   �  �  �            ��@@2    bb�     �B  l= �	   ��  �
     �   �   ���    $�   �  �  �            ���.�.2    kk�     &C  �? ;   ��  �
     �   �   ���    #�   �  �  �            ��tt2    t!t�     �C  B Ll   ��  �
     �   �   ���    "�   �  �  �            ����2    }(}�     "D  tD ��   ��  �
     �   �   ���    !�   �  �  �            ��'�'�2    �/�#�     �D  �F ��   ��  �
     �   �   ���     �   �  �  �            ���"*2    �@� �       =  Du  t�       M 
     J   �    C�#    � �   �  �  �             ��lc�2    �F� �       k  �v  �       M      J   �    C�#    � �   �  �  �             ��X��2    �L� �       �  x         M      J   �    C�$    � �   �  �  �             ���(�]2    �R� �       �  |y  L+       M      J   �    C�$    � �   �  �  �             ���:�2    �X� �       �  �z  �=       M      J   �    C�"    � �   �  �  �             ��l���2    �^� �       #  L|  �O       M      J   �    C�"    � �   �  �  �             ��U��2    �]� �       $  ��  z       N 
     K   �    �s�#    �   �  �  �             ����M2    �c� �       [  >�  d�       N      K   �    �s�#    �   �  �  �             ���i*�2    i� �       �  ċ  ��       N      K   �    �s�$    �   �  �  �             ��h��2    o� �       �  J�  �       N      K   �    �s�$    �   �  �  �             ���O�]2    u� �          Ў  `�       N      K   �    �s�"    �   �  �  �             ��1�3�2    {� �       7  V�  ��       N      K   �    �s�"    �   �  �  �             ���]�2    $�� �       �  ��  n=	       O 
     L   �    ��H#    � �   �  �  �             ��E�f�2    ,�� �       �  V�  
V	       O      L   �    ��H#    � �   �  �  �             ���$�72    4�� �       %  ��  �n	       O      L   �    ��H$    � �   �  �  �             ��%�!�2    <�� �       d  ��  B�	       O      L   �    ��H$    � �   �  �  �             ���*}2    D��       �  B�  ޟ	       O      L   �    ��H"    � �   �  �  �             ��	���2    L��       �  �  z�	       O      L   �    ��H"    � �   �  �  �             ����&2    R�      �  2�   C       P 
     M   �    ���#    �   �  �  �             ������2    Z�        ��  @_       P      M   �    ���#    �   �  �  �             ��b�U�2    b�      d  ��  `{       P      M   �    ���$    �   �  �  �             �����l2    j�       �  x�  ��       P      M   �    ���$    �   �  �  �             ��r!9�2    r�&      �  :�  ��       P      M   �    ���"    
�   �  �  �             �����[2    z�,       <  ��  ��       P      M   �    ���"    	�   �  �  �             ��=�4�2    �."n     �"  8�  ��       Q 
     N   �   ���#    �   �  �  �            ���F�&2    ��4(o     
#  �  ��       Q      N   �   ���#    �   �  �  �            ��%���2    ��:.p     \#  ��  x�       Q      N   �   ���$    �   �  �  �            ���|~+2    ��@4q     �#  ��  X�       Q      N   �   ���$    �   �  �  �            ��U	��2    ��F:r      $  ��  8       Q      N   �   ���"    �   �  �  �            ����	o52    ��L@s     R$  ��  /       Q      N   �   ���"    �   �  �  �            �����h2    ��MAx     Z)  ��  �'       R 
     O   �   �ؓ#    �   �  �  �            ��t,�2    ��SGy     �)  ��  �K       R      O   �   �ؓ#    �   �  �  �            �����V2    �YMz     *  ��  �o       R      O   �   �ؓ$    �   �  �  �            ���r	2�2    �_S{     k*  ��  \�       R      O   �   �ؓ$    �   �  �  �            ��M	
��2    �eY|     �*  ��  8�       R      O   �   �ؓ"    �   �  �  �            ���	�
='	2    �k_}     !+  ��  �       R      O   �   �ؓ"    �   �  �  �            ���kd2    �!l`�     �0  �  �       S 
     P      ���#    	�   �  �  �            ��>	��2    �)rf�     11  � �7       S      P      ���#    �   �  �  �            ����	Q"2    �1xl�     �1   
`       S      P      ���$    �   �  �  �            ���	�
��2    9~r�     �1  * �       S      P      ���$    �   �  �  �            ��J
=�|	2    A�x�     c2  F	 2�       S      P      ���"    �   �  �  �            ��"	&
2    I�~�     �2  b F�       S      P      ���"    �   �  �  �            ���C		�2    N���     9  n �L       T 
     Q   -   ���#    $�   �  �  �            ��	�	�a2    'V���     �9  �  y       T      Q   -   ���#    /�   �  �  �            ���	�
�2    0^���     �9  �! ��       T      Q   -   ���$    .�   �  �  �            ���
���	2    9f���     l:  $ 0�       T      Q   -   ���$    -�   �  �  �            ��[^e	t
2    Bn���     �:  V& ��       T      Q   -   ���"    ,�   �  �  �            ��&<
02    Kv���     P;  �( @+       T      Q   -   ���"    +�   �  �  �            ��W	'
��2    Qz���     CB  �; |�       U 
     R   .   ���#    �   �  �  �            ���	�
C.	2    Z����     �B  �= �       U      R   .   ���#    �   �  �  �            ���
���	2    c����     ?C  <@ �D       U      R   .   ���$    
�   �  �  �            �����	�
2    l����     �C  �B $v       U      R   .   ���$    	�   �  �  �            ��x�O
u2    u����     ;D  �D \�       U      R   .   ���"    �   �  �  �            ��X�B2    ~����     �D  DG ��       U      R   .   ���"    �   �  �  �            ��SX)
A2    ����     9  n �L       �

     �   �   ���#    %�   �  �  �            ��/G�
2    ����     �9  �  y       �
     �   �   ���#    $�   �  �  �            ��G��2    ���     �9  �! ��       �
     �   �   ���$    #�   �  �  �            ��a��2    ���     l:  $ 0�       �
     �   �   ���$    "�   �  �  �            ��t��2    �� �     �:  V& ��       �
     �   �   ���"    !�   �  �  �            ����2    ��'�     P;  �( @+       �
     �   �   ���"     �   �  �  �            ��X^/
G2    ����     CB  �; |�       �

        �   ���#    %�   �  �  �            ��6N�
2    ����     �B  �= �       �
        �   ���#    $�   �  �  �            ��"N��2    ���     ?C  <@ �D       �
        �   ���$    #�   �  �  �            ��h��2    ���     �C  �B $v       �
        �   ���$    "�   �  �  �            ��|��2    �� �     ;D  �D \�       �
        �   ���"    !�   �  �  �            ����2    ��'�     �D  DG ��       �
        �   ���"     �   �  �  �            ���8r2    � ��         Tt  D�       c 
     _   �    Cc#    � �   �  �  �             ��r[�2    � $��       N  �u  ��       c      _   �    Cc#    � �   �  �  �             ��C��2    � *��       }  $w  �       c      _   �    Cc$    � �   �  �  �             ����2    � 0��       �  �x         c      _   �    Cc$    � �   �  �  �             ���Mp�2    � 6��       �  �y  d1       c      _   �    Cc"    � �   �  �  �             ����[2    � <��       
  \{  �C       c      _   �    Cc"    � �   �  �  �             ���4N�2    	Z�       �    ^/	       e 
     a   �    �y #    � �   �  �  �             ����42    `'�       �  f�  �G	       e      a   �    �y #    � �   �  �  �             ��B��2    f/�         
�  �`	       e      a   �    �y $    � �   �  �  �             ���?�=2    l7�       @  ��  2y	       e      a   �    �y $    � �   �  �  �             �����2    !r?�         R�  Α	       e      a   �    �y "    � �   �  �  �             ��P�I2    'xG      �  ��  j�	       e      a   �    �y "    � �   �  �  �             ��0��2    )�M      �  B�   4       f 
     b   �    ��#    �   �  �  �             ��{m 2    /�U      �  �  @P       f      b   �    ��#    �   �  �  �             ���i�~2    5�]      >  ƶ  `l       f      b   �    ��$    �   �  �  �             ��9�*2    ;�e      �  ��  ��       f      b   �    ��$    �   �  �  �             ���O�2    A�m       �  J�  ��       f      b   �    ��"    
�   �  �  �             �����Y	2    G�u&        �  ��       f      b   �    ��"    	�   �  �  �             ���J�V2    I�z(n     �"  H�  �       g 
     c   �   ���#    �   �  �  �            ����7�2    O��.o     �"  (�  ��       g      c   �   ���#    �   �  �  �            ��W�f2    U��4p     3#  �  ��       g      c   �   ���$    �   �  �  �            ����j'	2    [��:q     �#  ��  h�       g      c   �   ���$    �   �  �  �            ��:	�	2    a��@r     �#  ��  H�       g      c   �   ���"    �   �  �  �            �����	{
2    g��Fs     )$  ��  (       g      c   �   ���"    �   �  �  �            ��/��22    h��Gx     0)  ��  �       h 
     d   �   ��X#    �   �  �  �            ���H�2    n��My     �)  ��  �:       h      d   �   ��X#    �   �  �  �            �����a	2    t��Sz     �)  ��  �^       h      d   �   ��X$    �   �  �  �            ��ySi	:
2    z��Y{     D*  ��  |�       h      d   �   ��X$    �   �  �  �            ����
�
2    ���_|     �*  ��  X�       h      d   �   ��X"    �   �  �  �            ��ic�
�2    ���e}     �*  ��  4�       h      d   �   ��X"    �   �  �  �            ���z^	2    ���f�     �0  ��  �       i 
     e      ���#    	�   �  �  �            ��$���	2    ���l�     1   &&       i      e      ���#    �   �  �  �            ���k�	m
2    � �r�     m1   :N       i      e      ���$    �   �  �  �            ��*q
]2    � x�     �1  : Nv       i      e      ���$    �   �  �  �            ����,)2    �	~�     ;2  V b�       i      e      ���"    �   �  �  �            ��3A	�2    ���     �2  r
 v�       i      e      ���"    �   �  �  �            ��N$>		
2    � ��     �8  ~ �9       j 
     f   /   ���#    $�   �  �  �            �����	�
2    �("��     X9  � `f       j      f   /   ���#    /�   �  �  �            ��8-�
}2    �0+��     �9  �  �       j      f   /   ���$    .�   �  �  �            ������2    �84��     <:  ,# p�       j      f   /   ���$    -�   �  �  �            ��k�	Wf2    �@=��     �:  f% ��       j      f   /   ���"    ,�   �  �  �            ��	4
4V2    �HF��      ;  �' �       j      f   /   ���"    +�   �  �  �            ����'
2    �NL��     B  �: ��       k 
     g   0   ���#    �   �  �  �            ��g[�
�2    �VU��     �B  �<         k      g   0   ���#    �   �  �  �            ������2    �^^��     C  L? <1       k      g   0   ���$    
�   �  �  �            ����	��2    �fg��     �C  �A tb       k      g   0   ���$    	�   �  �  �            ��=	m
��2    �np��     	D  �C ��       k      g   0   ���"    �   �  �  �            ���	(��2    vy��     �D  TF ��       k      g   0   ���"    �   �  �  �            ��	5
hy2    )����     �8  ~ �9       �

       �   ���#    %�   �  �  �            ���	�
X|2    0���     X9  � `f       �
       �   ���#    $�   �  �  �            ��f
�Y�2    7���     �9  �  �       �
       �   ���$    #�   �  �  �            ��V��2    >���     <:  ,# p�       �
       �   ���$    "�   �  �  �            ��!��S2    E���     �:  f% ��       �
       �   ���"    !�   �  �  �            ����(�2    L��!�      ;  �' �       �
       �   ���"     �   �  �  �            ��	9
n�2    )����     B  �: ��       �

       �   ���#    %�   �  �  �            ���	�
^�2    0���     �B  �<         �
       �   ���#    $�   �  �  �            ��k
�`�2    7���     C  L? <1       �
       �   ���$    #�   �  �  �            ��[��2    >���     �C  �A tb       �
       �   ���$    "�   �  �  �            ��'��]2    E���     	D  �C ��       �
       �   ���"    !�   �  �  �            �� �0�2    L��!�     �D  TF ��       �
       �   ���"     �   �  �  �             Q�Q�
2    �� ��       7  u  h�       } 
     w   �    ���    � �   �  �  �              ����
2    �� ��       f  pv  �       }      w   �    ���    � �   �  �  �              �1�1
2    �� ��       �  �w  �       }      w   �    ���    � �   �  �  �              $�$�
2    �� ��       �  @y  @(       }      w   �    ���    � �   �  �  �              n�n�
2    �� ��       �  �z  �:       }      w   �    ���    �    �  �  �              �;�;
2    �� ��       "  |  �L       }      w   �    ���    �   �  �  �              �-�-
2    �� ��         |�  �v       ~ 
     x   �    ���    �   �  �  �              xx
2    �� ��       S  �  �       ~      x   �    ���    �   �  �  �              U�U�
2    �� ��       �  ��  p�       ~      x   �    ���    �   �  �  �              �6�6
2    �� ��       �  �  Ķ       ~      x   �    ���    �   �  �  �              ��
2    �� ��       �  ��  �       ~      x   �    ���       �  �  �              h�h�
2    �� ��       /  �  l�       ~      x   �    ���      �  �  �              N�N�
2    �� ��       �  v�  �9	        
     y   �    ���    �   �  �  �              ��
2    �� ��       �  �  �R	             y   �    ���    �   �  �  �              �p�p
2    � ��         ��  "k	             y   �    ���    �   �  �  �              `�`�
2    ���       [  b�  ��	             y   �    ���    � 	  �  �  �              �X�X
2    �
��       �  �  Z�	             y   �    ���    � 
  �  �  �              '�'�
2    ��      �  ��  ��	             y   �    ���    �   �  �  �              �a�a
2    
      �  ��  `?       � 
     z   �    ���      �  �  �              /�/�
2            ��  �[       �      z   �    ���      �  �  �              �)�)
2    "      [  z�  �w       �      z   �    ���      �  �  �              ��
2    (       �  <�  ��       �      z   �    ���    	  �  �  �              x/x/
2    &.("      �  ��  �       �      z   �    ���    

  �  �  �              ����
2    .40(      3  ��   �       �      z   �    ���    	  �  �  �              oo
2    466*n     �"  ��  ��       � 
     {   �   ���      �  �  �             �s�s
2    <<>0o     �"  ��  ��       �      {   �   ���      �  �  �             9�9�
2    DBF6p     N#  ��  |�       �      {   �   ���      �  �  �             ����
2    LHN<q     �#  ��  \�       �      {   �   ���      �  �  �             BB
2    TNVBr     �#  |�  <       �      {   �   ���      �  �  �             ����
2    \T^Hs     A$  \�  +       �      {   �   ���      �  �  �             
�
�
2    aUcIx     Q)  ��  �#       � 
     |   �   ���      �  �  �             v1v1
2    i[kOy     �)  ��  lG       �      |   �   ���      �  �  �             ����
2    qasUz     	*  ��  Hk       �      |   �   ���      �  �  �             �c�c
2    yg{[{     e*  ��  $�       �      |   �   ���      �  �  �             ��
2    �m�a|     �*  ��   �       �      |   �   ���      �  �  �             ��	��	
2    �s�g}     +  ~�  ��       �      |   �   ���      �  �  �             �r�r
2    �t�h�     �0  �  n       � 
     }      ���    	  �  �  �             -�-�
2    �z�n�     (1  � �3       �      }      ���      �  �  �             ����
2    ���t�     �1  � �[       �      }      ���      �  �  �             ^J	^J	
2    ���z�     �1  � ��       �      }      ���      �  �  �             ��	��	
2    �����     ]2  
	 ��       �      }      ���      �  �  �             �	�
�	�

2    �����     �2  & ��       �      }      ���      �  �  �             b7b7
2    �����     
9  2 �G       � 
     ~   1   ���    $  �  �  �             ����
2    �����     |9  l pt       �      ~   1   ���    /  �  �  �             th	th	
2    �����     �9  �! ��       �      ~   1   ���    .  �  �  �             7	A
7	A

2    �����     `:  �# ��       �      ~   1   ���    -  �  �  �             �	�
�	�

2    �����     �:  & �       �      ~   1   ���    ,  �  �  �             �
��
�
2    �����     D;  T( �&       �      ~   1   ���    +  �  �  �             ��
2    �����     7B  P; ��       � 
        2   ���    $  �  �  �             ��	��	
2    ���     �B  �= �       �         2   ���    %  �  �  �             H	M
H	M

2    
���     3C   @  @       �         2   ���    
&  �  �  �             
:
:
2    ���     �C  XB 8q       �         2   ���    	'  �  �  �             �
�

2    ���     /D  �D p�       �         2   ���    (  �  �  �             ����
2    %�'��     �D  G ��       �         2   ���    )  �  �  �             �
��
�
2    WY �     
9  2 �G       �

       �   ���    %$  �  �  �             l�l�
2    `b�     |9  l pt       �
       �   ���    $%  �  �  �             9�9�
2    ik�     �9  �! ��       �
       �   ���    #&  �  �  �             R�R�
2    r!t�     `:  �# ��       �
       �   ���    "'  �  �  �             A�A�
2    {(}�     �:  & �       �
       �   ���    !(  �  �  �             @�@�
2    �/�#�     D;  T( �&       �
       �   ���     )  �  �  �             �
��
�
2    WY �     7B  P; ��       �

       �   ���    %$  �  �  �             r�r�
2    `b�     �B  �= �       �
       �   ���    $%  �  �  �             ?�?�
2    ik�     3C   @  @       �
       �   ���    #&  �  �  �             Y�Y�
2    r!t�     �C  XB 8q       �
       �   ���    "'  �  �  �             I�I�
2    {(}�     /D  �D p�       �
       �   ���    !(  �  �  �             I�I�
2    �/�#�     �D  G ��       �
       �   ���     )  �  �  �             �B�82    G�� �       F  �u  ��       � 
     �       ���    �    �  �  �             �r2    M�� �       u  �v  �	       �      �       ���    �    �  �  �             h�C�2    S�� �       �  Px         �      �       ���    �    �  �  �             �P�2    Y�� �       �  �y  X.       �      �       ���    �    �  �  �             $��M2    _�� �          {  �@       �      �       ���    �    �  �  �             ��2    e�� �       0  �|  �R       �      �       ���    �    �  �  �             n�I�2    m�� �       +  �  X}       � 
     �   	   ioe       �  �  �             �;��2    t�� �       a  z�  ��       �      �   	   ioe       �  �  �             ��A2    {�� �       �   �   �       �      �   	   ioe       �  �  �             ��2    ��� �       �  ��  T�       �      �   	   ioe       �  �  �             ��c�2    ��� �         �  ��       �      �   	   ioe       �  �  �             U��N2    ��� �       9  ��  ��       �      �   	   ioe       �  �  �             ��42    ��� �       �  �  �@	       � 
     �   
   ��    �    �  �  �             j��2    ��� �       �  ��  �Y	       �      �   
   ��    �    �  �  �             �dB�2    �� �       .  6�  *r	       �      �   
   ��    �    �  �  �             Q��?2    �� �       m  ڢ  Ɗ	       �      �   
   ��    �    �  �  �             �t��2    ��       �  ~�  b�	       �      �   
   ��    �    �  �  �             ;�P2    ��       �  "�  ��	       �      �   
   ��    �    �  �  �             �Q0�2    �$      �  n�  �F       � 
     �      :��       �  �  �             �{2    �,      &  0�   c       �      �      :��       �  �  �             �;�i2    �4      n  �          �      �      :��       �  �  �             #�9�2    �<       �  ��  @�       �      �      :��       �  �  �             �o�O2    �D&      �  v�  `�       �      �      :��    
   �  �  �             +	��2    �L,       F  8�  ��       �      �      :��    	   �  �  �             k�J2    �R."n     �"  t�  ��       � 
     �   �   ���       �  �  �             ����2    �Z4(o     #  T�  ��       �      �   �   ���       �  �  �             YW2    �b:.p     f#  4�  t�       �      �   �   ���       �  �  �             ���2    �j@4q     �#  �  T�       �      �   �   ���       �  �  �             �v	:2    �rF:r     
$  ��  4       �      �   �   ���       �  �  �             +	 
��2    �zL@s     \$  ��  3       �      �   �   ���       �  �  �             +�/�2    	MAx     f)   �   ,       � 
     �   �   ���       �  �  �             �s�H2    �SGy     �)  ��  �O       �      �   �   ���       �  �  �             5
	��2    �YMz     *  ��  �s       �      �   �   ���       �  �  �             ��	yS2    !�_S{     z*  ��  ��       �      �   �   ���       �  �  �             �	�
��2    )�eY|     �*  ��  p�       �      �   �   ���       �  �  �             >
Hic2    1�k_}     2+  ��  L�       �      �   �   ���       �  �  �             ���z2    5�l`�     �0   V       � 
     �      ���    	   �  �  �             �c	$�2    =�rf�     ?1  . j<       �      �      ���       �  �  �             	
�k2    E�xl�     �1  J ~d       �      �      ���       �  �  �             �	�
*2    M�~r�     2  f ��       �      �      ���       �  �  �             �
���2    U��x�     t2  �	 ��       �      �      ���       �  �  �             ]�3A	2    ]��~�     �2  � ��       �      �      ���       �  �  �             ��	N$2    a����     "9  � HQ       � 
     �   3   ���    $    �  �  �             e	V
��2    i����     �9  � �}       �      �   3   ���    /!   �  �  �             
8-2    q����     :  " X�       �      �   3   ���    ."   �  �  �             �
��2    y���     x:  X$ ��       �      �   3   ���    -#   �  �  �             ��k�	2    ����     �:  �& h       �      �   3   ���    ,$   �  �  �             ��	4
2    ����     \;  �( �/       �      �   3   ���    +%   �  �  �             �	�
��2    � ���     PB  �; h�       � 
     �   4   ���        �  �  �             Y
Wg[2    �)���     �B   > �       �      �   4   ���    !   �  �  �             "��2    �2���     LC  x@ �I       �      �   4   ���    
"   �  �  �             :��	2    �;���     �C  �B {       �      �   4   ���    	#   �  �  �             �'=	m
2    �D���     HD  (E H�       �      �   4   ���    $   �  �  �             �%�	(2    �M���     �D  �G ��       �      �   4   ���    %   �  �  �             ��	5
2    ���     "9  � HQ       �

       �   ���    %*   �  �  �             ���	�
2    ����     �9  � �}       �
       �   ���    $+   �  �  �             ��f
�2    ���     :  " X�       �
       �   ���    #,   �  �  �             �dV�2    ���     x:  X$ ��       �
       �   ���    "-   �  �  �             �!�2    �� �     �:  �& h       �
       �   ���    !.   �  �  �             O���2    �'�     \;  �( �/       �
       �   ���     /   �  �  �             ��	9
2    ���     PB  �; h�       �

       �   ���    %*   �  �  �             ���	�
2    ����     �B   > �       �
       �   ���    $+   �  �  �             ��k
�2    ���     LC  x@ �I       �
       �   ���    #,   �  �  �             l[�2    ���     �C  �B {       �
       �   ���    "-   �  �  �             $�'�2    �� �     HD  (E H�       �
       �   ���    !.   �  �  �             W� �2    �'�     �D  �G ��       �
       �   ���     /   �  �  �         ����   B D          O� r f       �  86  ��      
       ��            � .  �  �  �          ����   E G          V� v j       �  86  ��             ��            � /  �  �  �          ����   I J          ]� z n       �  86  ��             ��            � 0  �  �  �          ����   N P          d� ~ r       �  86  ��             ��            � 1  �  �  �          ����   R T          k� � v       �  86  ��             ��            � 2  �  �  �          ����   V X          r� � z       �  86  ��             ��            � 3  �  �  �          ����   H I          x� � u       �  �D  (�       
     	  ��	           	 � 8  �  �  �          ����   K M          � � y       �  �E  ��            	  ��	           	 � 9  �  �  �          ����   O P          �� � }         �F  @�            	  ��	           	 � :  �  �  �          ����   T V          �� � �       +  �G  ��            	  ��	           	 � ;  �  �  �          ����   Y Z          �� � �       F  �H  X�            	  ��	           	 � <  �  �  �          ����   ] _          �� � �       a  �I  ��            	  ��	           	 � =  �  �  �          ����   L M          �� � �       ,	  fS  b�   ��  
     
  ��           
 8  �  �  �         ����   O Q          � � �       M	  �T  F�   ��       
  ��           
 9  �  �  �         ����   S U          �� �       n	  �U  *�   ��       
  ��           
 :  �  �  �         ����   Y [          �� �       �	  �V  �   ��       
  ��           
 ;  �  �  �         ����   ^ _          �� �       �	  X  ��   ��       
  ��           
  <  �  �  �         ����   b d          �� �       �	  BY  ��   ��       
  ��           
 � =  �  �  �         ����   Q R          �� � n     �  �c  ��   ��   
       ���            B  �  �  �         ����   U V          �� � o     "  e   �   ��          ���            C  �  �  �         ����   Y [          �%� � p     J  bf  ��   ��          ���            D  �  �  �         ����   ` a          �+� � q     r  �g  �   ��          ���            
E  �  �  �         ����   d f          �1� � r     �  �h  ��   ��          ���            	F  �  �  �         ����   i k          �7� � s     �  @j   �   ��          ���            G  �  �  �         ����   U V          �7� � x     N  �u  ��   ��  !
       ���            B  �  �  y         ����   Y [          �=� � y     }  $w  �   ��  !       ���            C  �  �  y         ����   ^ _          C� � z     �  �x     ��  !       ���            D  �  �  y         ����   d f          I� � {     �  �y  d1   ��  !       ���            E  �  �  y         ����   i k          O� � |     
  \{  �C   ��  !       ���            F  �  �  y         ����   o p          U� � }     9  �|  �U   ��  !       ���            G  �  �  y         ����   Z \          &T� � �     5  0�  ��   ��  "
       ��'            "L  �  �  �         ����   _ `          .Z� � �     l  ��  ��   ��  "       ��'            !M  �  �  �         ����   d e          6`� � �     �  <�  H�   ��  "       ��'             N  �  �  �         ����   k l          >f� � �     �    ��   ��  "       ��'            O  �  �  �         ����   p r          Fl� � �       H�  ��   ��  "       ��'            P  �  �  �         ����   v w          Nr� � �     H  ΐ  D�   ��  "       ��'            Q  �  �  �         ����   _ `          U{� � �     �  *�  vD	   ��  #
       ��5            .L  �  �  �         ����   c e          ]�� � �     �  Ο  ]	   ��  #       ��5            -M  �  �  �         ����   h j          e�� � �     7  r�  �u	   ��  #       ��5            ,N  �  �  �         ����   o q          m�� � �     v  �  J�	   ��  #       ��5            +O  �  �  �         ����   u w          u�� �     �  ��  �	   ��  #       ��5            *P  �  �  �         ����   { }          }�� �     �  ^�  ��	   ��  #       ��5            )Q  �  �  �         ����   e g          ���     �  ��  �J   ��  $
       ��6            ;V  �  �  �         ����   j l          ���     0  l�  �f   ��  $       ��6            :W  �  �  �         ����   p q          ���     x  .�  ��   ��  $       ��6            9X  �  �  �         ����   w y          �� �     �  �   �   ��  $       ��6            8Y  �  �  �         ����   }           ��&�       ��   �   ��  $       ��6            7Z  �  �  �         ����   � �          ��, �     P  t�  @�   ��  $       ��6            6[  �  �  �         ����  A B          3� n b       �  D4  d�      �
       ��            � .  �  �  �          ����  D E          3� n b       �  D4  d�       �       ��            � /  �  �  �          ����  G I          3� n b       �  D4  d�   ��  �       ��            � 0  �  �  �          ����  L N          3� n b       �  D4  d�   ��  �       ��            � 1  �  �  �          ����  P R          3� n b       �  D4  d�   ��  �       ��            � 2  �  �  �          ����  T V          3� n b       �  D4  d�   ��  �       ��            � 3  �  �  �          ����  E F          c� � u       �  �B  ��   ��  �
     	  ��           	 � 8  �  �  �          ����  H J          j� � y       �  �C  ,�   ��  �     	  ��           	 � 9  �  �  �          ����  L M          q� � }       �  �D  ��   ��  �     	  ��           	 � :  �  �  �          ����  Q S          x� � �       �  �E  D�   ��  �     	  ��           	 � ;  �  �  �          ����  U W          � � �         �F  ��   ��  �     	  ��           	 � <  �  �  �          ����  Z [          �� � �       /  �G  \�   ��  �     	  ��           	 � =  �  �  �          ����  J L          �� � �       �  rQ  �   ��  �
     
  ��           
 8  �  �  �         ����  N O          � � �       	  �R  ʌ   ��  �     
  ��           
 9  �  �  �         ����  R S          �� �       7	  �S  ��   ��  �     
  ��           
 :  �  �  �         ����  X Y          �� �       X	  �T  ��   ��  �     
  ��           
 ;  �  �  �         ����  \ ^          �� �       y	  "V  v�   ��  �     
  ��           
  <  �  �  �         ����  a b          �� �       �	  NW  Z�   ��  �     
  ��           
 � =  �  �  �         ����  N P          �� � n     �  �a  8�   ��  �
       ���            B  �  �  �         ����  R T          �� � o     �  $c  ��   ��  �       ���            C  �  �  �         ����  V X          �%� � p       nd  (�   ��  �       ���            D  �  �  �         ����  \ ^          �+� � q     6  �e  ��   ��  �       ���            
E  �  �  �         ����  a c          �1� � r     ^  g  �   ��  �       ���            	F  �  �  �         ����  f h          �7� � s     �  Lh  ��   ��  �       ���            G  �  �  �         ����  T U          �7� � x       �s  (�   ��  �
       ���            B  �  �  {         ����  X Y          �=� � y     <  0u  p�   ��  �       ���            C  �  �  {         ����  \ ^          �C� � z     k  �v  �   ��  �       ���            D  �  �  {         ����  c d          �I� � {     �   x      ��  �       ���            E  �  �  {         ����  h i          O� � |     �  hy  H*   ��  �       ���            F  �  �  {         ����  m o          
U� � }     �  �z  �<   ��  �       ���            G  �  �  {         ����  X Y          T� � �     �  <�  He   ��  �
       ��,            "L  �  �  �         ����  \ ^          Z� � �     &    �z   ��  �       ��,            !M  �  �  �         ����  a b          !`� � �     ]  H�  ��   ��  �       ��,             N  �  �  �         ����  h i          )f� � �     �  ΋  D�   ��  �       ��,            O  �  �  �         ����  m n          1l� � �     �  T�  ��   ��  �       ��,            P  �  �  �         ����  r t          9r� � �       ڎ  ��   ��  �       ��,            Q  �  �  �         ����  ] _          @{� � �     n  6�  *'	   ��  �
       ��A            .L  �  �  �         ����  b c          H�� � �     �  ڝ  �?	   ��  �       ��A            -M  �  �  �         ����  g h          P�� � �     �  ~�  bX	   ��  �       ��A            ,N  �  �  �         ����  n o          X�� � �     +  "�  �p	   ��  �       ��A            +O  �  �  �         ����  s u          `�� �     j  Ƣ  ��	   ��  �       ��A            *P  �  �  �         ����  y {          h�� �     �  j�  6�	   ��  �       ��A            )Q  �  �  �         ����  c d          n��     �  ��  `+   ��  �
       ��B            ;V  �  �  �         ����  g i          v��     �  x�  �G   ��  �       ��B            :W  �  �  �         ����  m n          ~��     (  :�  �c   ��  �       ��B            9X  �  �  �         ����  t v          �� �     p  ��  �   ��  �       ��B            8Y  �  �  �         ����  z |          ��&�     �  ��  ��   ��  �       ��B            7Z  �  �  �         ����  � �          ��, �        ��   �   ��  �       ��B            6[  �  �  �         ����  B D          G� r f       �  �4  P�      �
       ��A            � .  �  �           ����  E G          N� v j       �  �5  ��       �       ��A            � /  �  �           ����  I J          U� z n       �  �6  0�   ��  �       ��A            � 0  �  �           ����  N P          \� ~ r         �7  ��   ��  �       ��A            � 1  �  �           ����  R T          c� � v         �8  �   ��  �       ��A            � 2  �  �           ����  V X          j� � z       /  �9  �   ��  �       ��A            � 3  �  �           ����  F H          p� � u       �  ,B  ��   ��  �
     	  ��B           	 � 8  �  �           ����  J K          w� � y       �  :C  D�   ��  �     	  ��B           	 � 9  �  �           ����  M O          ~� � }       �  HD  Ъ   ��  �     	  ��B           	 � :  �  �           ����  S T          �� � �       �  VE  \�   ��  �     	  ��B           	 � ;  �  �           ����  W Y          �� � �       
  dF  �   ��  �     	  ��B           	 � <  �  �           ����  [ ]          �� � �       %  rG  t�   ��  �     	  ��B           	 � =  �  �           ����  L M          �� � �       �  Q  �{   ��  �
     
  ��           
 8  �  �  �         ����  O Q          � � �       	  :R  ~�   ��  �     
  ��           
 9  �  �  �         ����  S U          �� �       ,	  fS  b�   ��  �     
  ��           
 :  �  �  �         ����  Y [          �� �       M	  �T  F�   ��  �     
  ��           
 ;  �  �  �         ����  ^ _          �� �       n	  �U  *�   ��  �     
  ��           
  <  �  �  �         ����  b d          �� �       �	  �V  �   ��  �     
  ��           
 � =  �  �  �         ����  P Q          �� � n     �  va  ��   ��  �
       ���            B  �  �  �         ����  T U          �� � o     �  �b   �   ��  �       ���            C  �  �  �         ����  X Y          �%� � p       
d  x�   ��  �       ���            D  �  �  �         ����  ^ `          �+� � q     *  Te  �   ��  �       ���            
E  �  �  �         ����  c d          �1� � r     R  �f  h�   ��  �       ���            	F  �  �  �         ����  h i          �7� � s     z  �g  ��   ��  �       ���            G  �  �  �         ����  U V          �7� � x        ds  �   ��  �
       ���            B  �  �  z         ����  Y [          �=� � y     /  �t  \�   ��  �       ���            C  �  �  z         ����  ^ _          �C� � z     ^  4v  �    ��  �       ���            D  �  �  z         ����  d f          I� � {     �  �w  �   ��  �       ���            E  �  �  z         ����  i k          O� � |     �  y  4%   ��  �       ���            F  �  �  z         ����  o p          U� � }     �  lz  |7   ��  �       ���            G  �  �  z         ����  Y Z          T� � �     �  ؆  �_   ��  �
       ��2            "L  �  �  �         ����  ^ _          &Z� � �       ^�  $u   ��  �       ��2            !M  �  �  �         ����  b d          .`� � �     O  �  x�   ��  �       ��2             N  �  �  �         ����  i k          6f� � �     �  j�  ̟   ��  �       ��2            O  �  �  �         ����  n p          >l� � �     �  ��   �   ��  �       ��2            P  �  �  �         ����  t v          Fr� � �     �  v�  t�   ��  �       ��2            Q  �  �  �         ����  _ `          M{� � �     _  қ  N!	   ��  �
       ��M            .L  �  �  �         ����  c e          U�� � �     �  v�  �9	   ��  �       ��M            -M  �  �  �         ����  h j          ]�� � �     �  �  �R	   ��  �       ��M            ,N  �  �  �         ����  o q          e�� � �       ��  "k	   ��  �       ��M            +O  �  �  �         ����  u w          m�� �     [  b�  ��	   ��  �       ��M            *P  �  �  �         ����  { }          u�� �     �  �  Z�	   ��  �       ��M            )Q  �  �  �         ����  d e          {��     �  R�   %   ��  �
       ��N            ;V  �  �  �         ����  i j          ���     �  �  @A   ��  �       ��N            :W  �  �  �         ����  n p          ���       ֵ  `]   ��  �       ��N            9X  �  �  �         ����  v w          �� �     `  ��  �y   ��  �       ��N            8Y  �  �  �         ����  | }          ��&�     �  Z�  ��   ��  �       ��N            7Z  �  �  �         ����  � �          ��, �     �  �  ��   ��  �       ��N            6[  �  �  �         ����  A B          5� r f       c  �;  �      ]
       ��T            � .  �  �            ����  D E          <� v j       y  �<  #       ]       ��T            � /  �  �            ����  G I          C� z n       �  �=  x+   ��  ]       ��T            � 0  �  �            ����  L N          J� ~ r       �  �>  �3   ��  ]       ��T            � 1  �  �            ����  P R          Q� � v       �  �?  X<   ��  ]       ��T            � 2  �  �            ����  T V          X� � z       �  �@  �D   ��  ]       ��T            � 3  �  �            ����  E F          ^� � u       R  4I  �   ��  ^
     	  ��U           	 � 8  �  �  !         ����  H J          e� � y       m  BJ  ��   ��  ^     	  ��U           	 � 9  �  �  !         ����  L M          l� � }       �  PK   �   ��  ^     	  ��U           	 � :  �  �  !         ����  Q S          s� � �       �  ^L  ��   ��  ^     	  ��U           	 � ;  �  �  !         ����  U W          z� � �       �  lM  8   ��  ^     	  ��U           	 � <  �  �  !         ����  Z [          �� � �       �  zN  �   ��  ^     	  ��U           	 � =  �  �  !         ����  J L          �� � �       �	  X  ��   ��  _
     
  ��           
 8  �  �  �         ����  N O          � � �       �	  BY  ��   ��  _     
  ��           
 9  �  �  �         ����  R S          �� �       �	  nZ  ��   ��  _     
  ��           
 :  �  �  �         ����  X Y          �� �       
  �[  ��   ��  _     
  ��           
 ;  �  �  �         ����  \ ^          �� �       4
  �\  ��   ��  _     
  ��           
  <  �  �  �         ����  a b          �� �       U
  �]  f	   ��  _     
  ��           
 � =  �  �  �         ����  N P          �� � n     �  ~h  ��   ��  `
       ���            B  �  �  �         ����  R T          �� � o     �  �i  `�   ��  `       ���            C  �  �  �         ����  V X          �%� � p     �  k  �   ��  `       ���            D  �  �  �         ����  \ ^          �+� � q       \l  P   ��  `       ���            
E  �  �  �         ����  a c          �1� � r     *  �m  �#   ��  `       ���            	F  �  �  �         ����  f h          �7� � s     R  �n  @3   ��  `       ���            G  �  �  �         ����  T U          �7� � x     �  lz  |7   ��  a
       ���            B  �  �  |         ����  X Y          �=� � y       �{  �I   ��  a       ���            C  �  �  |         ����  \ ^          �C� � z     H  <}  \   ��  a       ���            D  �  �  |         ����  c d          �I� � {     w  �~  Tn   ��  a       ���            E  �  �  |         ����  h i          �O� � |     �  �  ��   ��  a       ���            F  �  �  |         ����  m o          U� � }     �  t�  �   ��  a       ���            G  �  �  |         ����  X Y          T� � �     �  ��  @�   ��  b
       ��7            "L  �  �  �         ����  \ ^          Z� � �       f�  ��   ��  b       ��7            !M  �  �  �         ����  a b          `� � �     K  �  ��   ��  b       ��7             N  �  �  �         ����  h i          $f� � �     �  r�  <   ��  b       ��7            O  �  �  �         ����  m n          ,l� � �     �  ��  �   ��  b       ��7            P  �  �  �         ����  r t          4r� � �     �  ~�  �,   ��  b       ��7            Q  �  �  �         ����  ] _          ;{� � �     m  ڢ  Ɗ	   ��  c
       ��Y            .L  �  �  �         ����  b c          C�� � �     �  ~�  b�	   ��  c       ��Y            -M  �  �  �         ����  g h          K�� � �     �  "�  ��	   ��  c       ��Y            ,N  �  �  �         ����  n o          S�� � �     *  Ƨ  ��	   ��  c       ��Y            +O  �  �  �         ����  s u          [�� �     i  j�  6�	   ��  c       ��Y            *P  �  �  �         ����  y {          c�� �     �  �  �
   ��  c       ��Y            )Q  �  �  �         ����  c d          i��     �  Z�  ��   ��  d
       ��Z            ;V  �  �  �         ����  g i          q��     �  �  ��   ��  d       ��Z            :W  �  �  �         ����  m n          y��     8  ޼  ��   ��  d       ��Z            9X  �  �  �         ����  t v          �� �     �  ��   �   ��  d       ��Z            8Y  �  �  �         ����  z |          ��&�     �  b�      ��  d       ��Z            7Z  �  �  �         ����  � �          ��, �       $�  @"   ��  d       ��Z            6[  �  �  �         ����  D E          U� n b       )  X9        �
       ��g            � .  �  �  3         ����  G H          U� n b       )  X9        �       ��g            � /  �  �  3         ����  J L          U� n b       )  X9        �       ��g            � 0  �  �  3         ����  P Q          U� n b       )  X9        �       ��g            � 1  �  �  3         ����  T U          U� n b       )  X9        �       ��g            � 2  �  �  3         ����  X Z          U� n b       )  X9        �       ��g            � 3  �  �  3         ����  I J          �� � u       *  �G  h�   ��  �
       ��h           	 � 8  �  �  4         ����  M N          �� � y       E  �H  ��   ��  �       ��h           	 � 9  �  �  4         ����  P R          �� � }       `  �I  ��   ��  �       ��h           	 � :  �  �  4         ����  V X          �� � �       {  �J  �   ��  �       ��h           	 � ;  �  �  4         ����  Z \          �� � �       �  �K  ��   ��  �       ��h           	 � <  �  �  4         ����  _ a          �� � �       �  �L  $   ��  �       ��h           	 � =  �  �  4         ����  M N          �� � �       �	  �V  ·   ��  �
     	  ��           
 8  �  �           ����  Q R          � � �       �	  �W  ��   ��  �     	  ��           
 9  �  �           ����  U V          �� �       �	  �X  ��   ��  �     	  ��           
 :  �  �           ����  [ \          �� �       �	  
Z  n�   ��  �     	  ��           
 ;  �  �           ����  _ a          �� �       
  6[  R�   ��  �     	  ��           
  <  �  �           ����  d f          �� �       )
  b\  6�   ��  �     	  ��           
 � =  �  �           ����  R T          �� � n     Z  �f  (�   ��  �
     
  ���            B  �  �  �         ����  V X          �� � o     �  8h  ��   ��  �     
  ���            C  �  �  �         ����  [ \          �%� � p     �  �i  �   ��  �     
  ���            D  �  �  �         ����  a c          �+� � q     �  �j  �   ��  �     
  ���            
E  �  �  �         ����  f h          �1� � r     �  l     ��  �     
  ���            	F  �  �  �         ����  k m          �7� � s     "  `m  �    ��  �     
  ���            G  �  �  �         ����  V X          7� � x     �  �x  ,#   ��  �
       ���            B  �  �  ~         ����  [ \          =� � y     �  Dz  t5   ��  �       ���            C  �  �  ~         ����  _ a          C� � z       �{  �G   ��  �       ���            D  �  �  ~         ����  f h          I� � {     C  }  Z   ��  �       ���            E  �  �  ~         ����  k m          $O� � |     r  |~  Ll   ��  �       ���            F  �  �  ~         ����  p r          ,U� � }     �  �  �~   ��  �       ���            G  �  �  ~         ����  \ ]          3T� � �     �  P�  `�   ��  �
       ��<            "L  �  �  �         ����  ` b          ;Z� � �     �  ֍  ��   ��  �       ��<            !M  �  �  �         ����  e g          C`� � �       \�  �   ��  �       ��<             N  �  �  �         ����  l n          Kf� � �     J  �  \�   ��  �       ��<            O  �  �  �         ����  r s          Sl� � �     �  h�  �   ��  �       ��<            P  �  �  �         ����  w y          [r� � �     �  �     ��  �       ��<            Q  �  �  �         ����  ` a          b{� � �     1  J�  Vs	   ��  �
       ��e            .L  �  �  �         ����  e f          j�� � �     p  �  �	   ��  �       ��e            -M  �  �  �         ����  j k          r�� � �     �  ��  ��	   ��  �       ��e            ,N  �  �  �         ����  q s          z�� � �     �  6�  *�	   ��  �       ��e            +O  �  �  �         ����  w x          ��� �     -  ڧ  ��	   ��  �       ��e            *P  �  �  �         ����  } ~          ��� �     l  ~�  b�	   ��  �       ��e            )Q  �  �  �         ����  g h          ���     h  ʷ  �|   ��  �
       ��f            ;V  �  �  �         ����  l m          ���     �  ��  ��   ��  �       ��f            :W  �  �  �         ����  q s          ���     �  N�  �   ��  �       ��f            9X  �  �  �         ����  y {          �� �     @  �   �   ��  �       ��f            8Y  �  �  �         ����   �          ��&�     �  Ҿ   �   ��  �       ��f            7Z  �  �  �         ����  � �          ��, �     �  ��  @	   ��  �       ��f            6[  �  �  �         ����  B D          ;� n b         �7  �      )
       ��z            � .  �  �  F         ����  E G          ;� n b         �7  �      )       ��z            � /  �  �  F         ����  I J          ;� n b         �7  �      )       ��z            � 0  �  �  F         ����  N P          ;� n b         �7  �      )       ��z            � 1  �  �  F         ����  R T          ;� n b         �7  �      )       ��z            � 2  �  �  F         ����  V X          ;� n b         �7  �      )       ��z            � 3  �  �  F         ����  F H          k� � u         F  ȼ   ��  *
     	  ��{           	 � 8  �  �  G         ����  J K          r� � y         "G  T�   ��  *     	  ��{           	 � 9  �  �  G         ����  M O          y� � }       8  0H  ��   ��  *     	  ��{           	 � :  �  �  G         ����  S T          �� � �       S  >I  l�   ��  *     	  ��{           	 � ;  �  �  G         ����  W Y          �� � �       n  LJ  ��   ��  *     	  ��{           	 � <  �  �  G         ����  [ ]          �� � �       �  ZK  ��   ��  *     	  ��{           	 � =  �  �  G         ����  L M          �� � �       X	  �T  ��   ��  +
     
  ��           
 8  �  �  
         ����  O Q          � � �       y	  "V  v�   ��  +     
  ��           
 9  �  �  
         ����  S U          �� �       �	  NW  Z�   ��  +     
  ��           
 :  �  �  
         ����  Y [          �� �       �	  zX  >�   ��  +     
  ��           
 ;  �  �  
         ����  ^ _          �� �       �	  �Y  "�   ��  +     
  ��           
  <  �  �  
         ����  b d          �� �       �	  �Z  �   ��  +     
  ��           
 � =  �  �  
         ����  P Q          �� � n     *  ^e  h�   ��  ,
       ���            B  �  �  �         ����  T U          �� � o     R  �f  ��   ��  ,       ���            C  �  �  �         ����  X Y          �%� � p     z  �g  X�   ��  ,       ���            D  �  �  �         ����  ^ `          �+� � q     �  <i  ��   ��  ,       ���            
E  �  �  �         ����  c d          �1� � r     �  �j  H�   ��  ,       ���            	F  �  �  �         ����  h i          �7� � s     �  �k  �   ��  ,       ���            G  �  �  �         ����  U V          �7� � x     �  Lw  �   ��  -
       ���            B  �  �  }         ����  Y [          �=� � y     �  �x  $!   ��  -       ���            C  �  �  }         ����  ^ _          �C� � z     �  z  l3   ��  -       ���            D  �  �  }         ����  d f          I� � {       �{  �E   ��  -       ���            E  �  �  }         ����  i k          
O� � |     >  �|  �W   ��  -       ���            F  �  �  }         ����  o p          U� � }     m  T~  Dj   ��  -       ���            G  �  �  }         ����  Y Z          T� � �     m  ��  ��   ��  .
       ��A            "L  �  �  �         ����  ^ _          !Z� � �     �  F�  ԫ   ��  .       ��A            !M  �  �  �         ����  b d          )`� � �     �  ̍  (�   ��  .       ��A             N  �  �  �         ����  i k          1f� � �       R�  |�   ��  .       ��A            O  �  �  �         ����  n p          9l� � �     I  ؐ  ��   ��  .       ��A            P  �  �  �         ����  t v          Ar� � �     �  ^�  $   ��  .       ��A            Q  �  �  �         ����  _ `          H{� � �     �  ��  �[	   ��  /
       ��q            .L  �  �           ����  c e          P�� � �     4  ^�  �t	   ��  /       ��q            -M  �  �           ����  h j          X�� � �     s  �  �	   ��  /       ��q            ,N  �  �           ����  o q          `�� � �     �  ��  ��	   ��  /       ��q            +O  �  �           ����  u w          h�� �     �  J�  V�	   ��  /       ��q            *P  �  �           ����  { }          p�� �     0  �  ��	   ��  /       ��q            )Q  �  �           ����  d e          v��     (  :�  �c   ��  0
       ��r            ;V  �  �           ����  i j          ~��     p  ��  �   ��  0       ��r            :W  �  �           ����  n p          ���     �  ��  ��   ��  0       ��r            9X  �  �           ����  v w          �� �        ��   �   ��  0       ��r            8Y  �  �           ����  | }          ��&�     H  B�   �   ��  0       ��r            7Z  �  �           ����  � �          ��, �     �  �  @�   ��  0       ��r            6[  �  �           ����  B D          M� n b       q  x<  8       �
     �   �            � .  �  �  Y         ����  E G          M� n b       q  x<  8       �     �   �            � /  �  �  Y         ����  I J          M� n b       q  x<  8       �     �   �            � 0  �  �  Y         ����  N P          M� n b       q  x<  8       �     �   �            � 1  �  �  Y         ����  R T          M� n b       q  x<  8       �     �   �            � 2  �  �  Y         ����  V X          M� n b       q  x<  8       �     �   �            � 3  �  �  Y         ����  H I          }� � u       z  �J  ��   ��  �
     �   �           	 � 8  �  �  Z         ����  K M          �� � y       �  �K  4�   ��  �     �   �           	 � 9  �  �  Z         ����  O P          �� � }       �  �L  �    ��  �     �   �           	 � :  �  �  Z         ����  T V          �� � �       �  �M  L   ��  �     �   �           	 � ;  �  �  Z         ����  Y Z          �� � �       �  �N  �   ��  �     �   �           	 � <  �  �  Z         ����  ] _          �� � �         
P  d    ��  �     �   �           	 � =  �  �  Z         ����  L M          �� � �       �	  �Y  "�   ��  �
     �   �           
 8  �  �  �         ����  O Q          � � �       �	  �Z  �   ��  �     �   �           
 9  �  �  �         ����  S U          �� �       
  �[  ��   ��  �     �   �           
 :  �  �  �         ����  Y [          �� �       ?
  *]  �    ��  �     �   �           
 ;  �  �  �         ����  ^ _          �� �       `
  V^  �   ��  �     �   �           
  <  �  �  �         ����  b d          �� �       �
  �_  �   ��  �     �   �           
 � =  �  �  �         ����  Q R          �� � n     �  j  ��   ��  �
     �   �            B  �  �  �         ����  U V          �� � o     �  Xk      ��  �     �   �            C  �  �  �         ����  Y [          �%� � p     
  �l  �   ��  �     �   �            D  �  �  �         ����  ` a          �+� � q     2  �m  '   ��  �     �   �            
E  �  �  �         ����  d f          �1� � r     Z  6o  �6   ��  �     �   �            	F  �  �  �         ����  i k          �7� � s     �  �p   F   ��  �     �   �            G  �  �  �         ����  U V          �7� � x       �{  �K   ��  �
     �   �            B  �  �           ����  Y [          =� � y     M  d}  ^   ��  �     �   �            C  �  �           ����  ^ _          C� � z     |  �~  \p   ��  �     �   �            D  �  �           ����  d f          I� � {     �  4�  ��   ��  �     �   �            E  �  �           ����  i k          O� � |     �  ��  �   ��  �     �   �            F  �  �           ����  o p          $U� � }     	  �  4�   ��  �     �   �            G  �  �           ����  Z \          +T� � �       p�   �   ��  �
     �   F            "L  �  �  �         ����  _ `          3Z� � �     L  ��  t�   ��  �     �   F            !M  �  �  �         ����  d e          ;`� � �     �  |�  �   ��  �     �   F             N  �  �  �         ����  k l          Cf� � �     �  �     ��  �     �   F            O  �  �  �         ����  p r          Kl� � �     �  ��  p-   ��  �     �   F            P  �  �  �         ����  v w          Sr� � �     (  �  �B   ��  �     �   F            Q  �  �  �         ����  _ `          Z{� � �     �  j�  6�	   ��  �
     �   }            .L  �  �           ����  c e          b�� � �     �  �  Һ	   ��  �     �   }            -M  �  �           ����  h j          j�� � �     '  ��  n�	   ��  �     �   }            ,N  �  �           ����  o q          r�� � �     f  V�  
�	   ��  �     �   }            +O  �  �           ����  u w          z�� �     �  ��  �
   ��  �     �   }            *P  �  �           ����  { }          ��� �     �  ��  B
   ��  �     �   }            )Q  �  �           ����  e g          ���     �  �  ��   ��  �
     �   ~            ;V  �  �           ����  j l          ���     0  ��  ��   ��  �     �   ~            :W  �  �           ����  p q          ���     x  n�  ��   ��  �     �   ~            9X  �  �           ����  w y          �� �     �  0�      ��  �     �   ~            8Y  �  �           ����  }           ��&�       ��      ��  �     �   ~            7Z  �  �           ����  � �          ��, �     P  ��  @;   ��  �     �   ~            6[  �  �           ����   9 :          � � Hl       �  (7  h�      1
       ��            � .  �  �  �          ����   < =          � � Op         8  ��       1       ��            � /  �  �  �          ����   ? @          � � Vt       #  9  H   ��  1       ��            � 0  �  �  �          ����   C D          � � ]x       9  �9  �	   ��  1       ��            � 1  �  �  �          ����   F H          � � d|       O  �:  (   ��  1       ��            � 2  �  �  �          ����   J K          � � k�       e  �;  �   ��  1       ��            � 3  �  �  �          ����   = >          � � q{       �  �D  (�   ��  2
     	  ��           	 � 8  �  �  �          ����   @ A          � � x       �  �E  ��   ��  2     	  ��           	 � 9  �  �  �          ����   C D          � � �         �F  @�   ��  2     	  ��           	 � :  �  �  �          ����   H I          � � ��       +  �G  ��   ��  2     	  ��           	 � ;  �  �  �          ����   K M          � � ��       F  �H  X�   ��  2     	  ��           	 � <  �  �  �          ����   O Q          � � ��       a  �I  ��   ��  2     	  ��           	 � =  �  �  �          ����   A B          � � ��       ,	  fS  b�   ��  3
     
  ��           
 8  �  �  �         ����   D E          � � ��       M	  �T  F�   ��  3     
  ��           
 9  �  �  �         ����   G I          � � ��       n	  �U  *�   ��  3     
  ��           
 :  �  �  �         ����   L N          � ��       �	  �V  �   ��  3     
  ��           
 ;  �  �  �         ����   P R          � ��       �	  X  ��   ��  3     
  ��           
  <  �  �  �         ����   T V          � ��       �	  BY  ��   ��  3     
  ��           
 � =  �  �  �         ����   E F          � �� n     �  �c  ��   ��  4
       ���            B  �  �  �         ����   H J          � �� o     "  e   �   ��  4       ���            C  �  �  �         ����   L M          �  �� p     J  bf  ��   ��  4       ���            D  �  �  �         ����   Q S          � &�� q     r  �g  �   ��  4       ���            
E  �  �  �         ����   U W          � ,�� r     �  �h  ��   ��  4       ���            	F  �  �  �         ����   Z [          � 2�� s     �  @j   �   ��  4       ���            G  �  �  �         ����   I J          � 3�� x     N  �u  ��   ��  5
       ���            B  �  �  �         ����   M N          � 9�� y     }  $w  �   ��  5       ���            C  �  �  �         ����   P R          � ? � z     �  �x     ��  5       ���            D  �  �  �         ����   V X          � E� {     �  �y  d1   ��  5       ���            E  �  �  �         ����   Z \          � K� |     
  \{  �C   ��  5       ���            F  �  �  �         ����   _ a          Q� }     9  �|  �U   ��  5       ���            G  �  �  �         ����   L M          � Q� �     5  0�  ��   ��  6
       ��(            "L  �  �  �         ����   O Q          W'� �     l  ��  ��   ��  6       ��(            !M  �  �  �         ����   S U          	]/� �     �  <�  H�   ��  6       ��(             N  �  �  �         ����   Y [          c7� �     �    ��   ��  6       ��(            O  �  �  �         ����   ^ _          i?� �       H�  ��   ��  6       ��(            P  �  �  �         ����   b d          oG� �     H  ΐ  D�   ��  6       ��(            Q  �  �  �         ����   Q R           oN� �     �  *�  vD	   ��  7
       ��7            .L  �  �  �         ����   U V          &uV� �     �  Ο  ]	   ��  7       ��7            -M  �  �  �         ����   Y [          ,{^� �     7  r�  �u	   ��  7       ��7            ,N  �  �  �         ����   ` a          2�f� �     v  �  J�	   ��  7       ��7            +O  �  �  �         ����   d f          8�n� �     �  ��  �	   ��  7       ��7            *P  �  �  �         ����   i k          >�v�     �  ^�  ��	   ��  7       ��7            )Q  �  �  �         ����   U V          @�|�     �  ��  �J   ��  8
       ��8            ;V  �  �  �         ����   Y [          F���     0  l�  �f   ��  8       ��8            :W  �  �  �         ����   ^ _          L���     x  .�  ��   ��  8       ��8            9X  �  �  �         ����   d f          R���     �  �   �   ��  8       ��8            8Y  �  �  �         ����   i k          X�� �       ��   �   ��  8       ��8            7Z  �  �  �         ����   o p          ^��&�     P  t�  @�   ��  8       ��8            6[  �  �  �         ����  9 :          { � 3l       �  45  ��      �
       ��             � .  �  �  �          ����  < =           � :p       �  $6  D�       �       ��             � /  �  �  �          ����  ? @          � � At       �  7  ��   ��  �       ��             � 0  �  �  �          ����  C D          � � Hx         8  $�   ��  �       ��             � 1  �  �  �          ����  F H          � � O|       "  �8  �    ��  �       ��             � 2  �  �  �          ����  J K          � � V�       8  �9  	   ��  �       ��             � 3  �  �  �          ����  = >          � � \{       �  �B  ��   ��  �
     	  ��!           	 � 8  �  �  �          ����  @ A          � � c       �  �C  ,�   ��  �     	  ��!           	 � 9  �  �  �          ����  C D          � � j�       �  �D  ��   ��  �     	  ��!           	 � :  �  �  �          ����  H I          � � q�       �  �E  D�   ��  �     	  ��!           	 � ;  �  �  �          ����  K M          � � x�         �F  ��   ��  �     	  ��!           	 � <  �  �  �          ����  O Q          � � �       /  �G  \�   ��  �     	  ��!           	 � =  �  �  �          ����  ? A          � � ��       �  rQ  �   ��  �
     
  ��	           
 8  �  �  �         ����  C D          � � ��       	  �R  ʌ   ��  �     
  ��	           
 9  �  �  �         ����  F G          � � ��       7	  �S  ��   ��  �     
  ��	           
 :  �  �  �         ����  K L          � � ��       X	  �T  ��   ��  �     
  ��	           
 ;  �  �  �         ����  O P          � � ��       y	  "V  v�   ��  �     
  ��	           
  <  �  �  �         ����  S T          � � ��       �	  NW  Z�   ��  �     
  ��	           
 � =  �  �  �         ����  D E          � � �� n     �  �a  8�   ��  �
       ���            B  �  �  �         ����  G H          � �� o     �  $c  ��   ��  �       ���            C  �  �  �         ����  J L          � �� p       nd  (�   ��  �       ���            D  �  �  �         ����  P Q          � �� q     6  �e  ��   ��  �       ���            
E  �  �  �         ����  T U          � �� r     ^  g  �   ��  �       ���            	F  �  �  �         ����  X Z          � �� s     �  Lh  ��   ��  �       ���            G  �  �  �         ����  H I          � �� x       �s  (�   ��  �
       ���            B  �  �  �         ����  K M          � $�� y     <  0u  p�   ��  �       ���            C  �  �  �         ����  O P          � *�� z     k  �v  �   ��  �       ���            D  �  �  �         ����  T V          � 0�� {     �   x      ��  �       ���            E  �  �  �         ����  Y Z          � 6�� |     �  hy  H*   ��  �       ���            F  �  �  �         ����  ] _          � <� }     �  �z  �<   ��  �       ���            G  �  �  �         ����  L M          � <
� �     �  <�  He   ��  �
       ��-            "L  �  �  �         ����  O Q          � B� �     &    �z   ��  �       ��-            !M  �  �  �         ����  S U          � H� �     ]  H�  ��   ��  �       ��-             N  �  �  �         ����  Y [          � N"� �     �  ΋  D�   ��  �       ��-            O  �  �  �         ����  ^ _          � T*� �     �  T�  ��   ��  �       ��-            P  �  �  �         ����  b d          Z2� �       ڎ  ��   ��  �       ��-            Q  �  �  �         ����  Q R          Z9� �     n  6�  *'	   ��  �
       ��C            .L  �  �  �         ����  U V          `A� �     �  ڝ  �?	   ��  �       ��C            -M  �  �  �         ����  Y [          fI� �     �  ~�  bX	   ��  �       ��C            ,N  �  �  �         ����  ` a          lQ� �     +  "�  �p	   ��  �       ��C            +O  �  �  �         ����  d f          #rY� �     j  Ƣ  ��	   ��  �       ��C            *P  �  �  �         ����  i k          )xa�     �  j�  6�	   ��  �       ��C            )Q  �  �  �         ����  T U          +�g�     �  ��  `+   ��  �
       ��D            ;V  �  �  �         ����  X Y          1�o�     �  x�  �G   ��  �       ��D            :W  �  �  �         ����  \ ^          7�w�     (  :�  �c   ��  �       ��D            9X  �  �  �         ����  c d          =��     p  ��  �   ��  �       ��D            8Y  �  �  �         ����  h i          C�� �     �  ��  ��   ��  �       ��D            7Z  �  �  �         ����  m o          I��&�        ��   �   ��  �       ��D            6[  �  �  �         ����  9 :          � � @l       �  �4  P�      
       ��F            � .  �  �           ����  < =          � � Gp       �  �5  ��              ��F            � /  �  �           ����  ? @          � � Nt       �  �6  0�   ��         ��F            � 0  �  �           ����  C D          � � Ux         �7  ��   ��         ��F            � 1  �  �           ����  F H          � � \|         �8  �   ��         ��F            � 2  �  �           ����  J K          � � c�       /  �9  �   ��         ��F            � 3  �  �           ����  = >          � � i{       �  ,B  ��   ��  	
     	  ��G           	 � 8  �  �           ����  @ A          � � p       �  :C  D�   ��  	     	  ��G           	 � 9  �  �           ����  C D          � � w�       �  HD  Ъ   ��  	     	  ��G           	 � :  �  �           ����  H I          � � ~�       �  VE  \�   ��  	     	  ��G           	 � ;  �  �           ����  K M          � � ��       
  dF  �   ��  	     	  ��G           	 � <  �  �           ����  O Q          � � ��       %  rG  t�   ��  	     	  ��G           	 � =  �  �           ����  ? A          � � ��       �  Q  �{   ��  

     
  ��           
 8  �  �  �         ����  C D          � � ��       	  :R  ~�   ��  
     
  ��           
 9  �  �  �         ����  F G          � � ��       ,	  fS  b�   ��  
     
  ��           
 :  �  �  �         ����  K L          � � ��       M	  �T  F�   ��  
     
  ��           
 ;  �  �  �         ����  O P          �  ��       n	  �U  *�   ��  
     
  ��           
  <  �  �  �         ����  S T          � ��       �	  �V  �   ��  
     
  ��           
 � =  �  �  �         ����  D E          � �� n     �  va  ��   ��  
       ���            B  �  �  �         ����  G H          � �� o     �  �b   �   ��         ���            C  �  �  �         ����  J L          � �� p       
d  x�   ��         ���            D  �  �  �         ����  P Q          � �� q     *  Te  �   ��         ���            
E  �  �  �         ����  T U          � $�� r     R  �f  h�   ��         ���            	F  �  �  �         ����  X Z          � *�� s     z  �g  ��   ��         ���            G  �  �  �         ����  H I          � +�� x        ds  �   ��  
       ���            B  �  �  �         ����  K M          � 1�� y     /  �t  \�   ��         ���            C  �  �  �         ����  O P          � 7�� z     ^  4v  �    ��         ���            D  �  �  �         ����  T V          � = � {     �  �w  �   ��         ���            E  �  �  �         ����  Y Z          � C� |     �  y  4%   ��         ���            F  �  �  �         ����  ] _          � I� }     �  lz  |7   ��         ���            G  �  �  �         ����  L M          � I� �     �  ؆  �_   ��  
       ��3            "L  �  �  �         ����  O Q          � O� �       ^�  $u   ��         ��3            !M  �  �  �         ����  S U          U'� �     O  �  x�   ��         ��3             N  �  �  �         ����  Y [          [/� �     �  j�  ̟   ��         ��3            O  �  �  �         ����  ^ _          a7� �     �  ��   �   ��         ��3            P  �  �  �         ����  b d          g?� �     �  v�  t�   ��         ��3            Q  �  �  �         ����  Q R          gF� �     _  қ  N!	   ��  
       ��O            .L  �  �  �         ����  U V          mN� �     �  v�  �9	   ��         ��O            -M  �  �  �         ����  Y [          $sV� �     �  �  �R	   ��         ��O            ,N  �  �  �         ����  ` a          *y^� �       ��  "k	   ��         ��O            +O  �  �  �         ����  d f          0f� �     [  b�  ��	   ��         ��O            *P  �  �  �         ����  i k          6�n�     �  �  Z�	   ��         ��O            )Q  �  �  �         ����  T U          8�t�     �  R�   %   ��  
       ��P            ;V  �  �  �         ����  X Y          >�|�     �  �  @A   ��         ��P            :W  �  �  �         ����  \ ^          D���       ֵ  `]   ��         ��P            9X  �  �  �         ����  c d          J���     `  ��  �y   ��         ��P            8Y  �  �  �         ����  h i          P�� �     �  Z�  ��   ��         ��P            7Z  �  �  �         ����  m o          V��&�     �  �  ��   ��         ��P            6[  �  �  �         ����  9 :          v � .l       c  �;  �      n
       ��Y            � .  �  �  %         ����  < =          z � 5p       y  �<  #       n       ��Y            � /  �  �  %         ����  ? @          ~ � <t       �  �=  x+   ��  n       ��Y            � 0  �  �  %         ����  C D          � � Cx       �  �>  �3   ��  n       ��Y            � 1  �  �  %         ����  F H          � � J|       �  �?  X<   ��  n       ��Y            � 2  �  �  %         ����  J K          � � Q�       �  �@  �D   ��  n       ��Y            � 3  �  �  %         ����  = >          � � W{       R  4I  �   ��  o
     	  ��Z           	 � 8  �  �  &         ����  @ A          � � ^       m  BJ  ��   ��  o     	  ��Z           	 � 9  �  �  &         ����  C D          � � e�       �  PK   �   ��  o     	  ��Z           	 � :  �  �  &         ����  H I          � � l�       �  ^L  ��   ��  o     	  ��Z           	 � ;  �  �  &         ����  K M          � � s�       �  lM  8   ��  o     	  ��Z           	 � <  �  �  &         ����  O Q          � � z�       �  zN  �   ��  o     	  ��Z           	 � =  �  �  &         ����  ? A          � � �       �	  X  ��   ��  p
     
  ��           
 8  �  �            ����  C D          � � ��       �	  BY  ��   ��  p     
  ��           
 9  �  �            ����  F G          � � ��       �	  nZ  ��   ��  p     
  ��           
 :  �  �            ����  K L          � � ��       
  �[  ��   ��  p     
  ��           
 ;  �  �            ����  O P          � � ��       4
  �\  ��   ��  p     
  ��           
  <  �  �            ����  S T          � � ��       U
  �]  f	   ��  p     
  ��           
 � =  �  �            ����  D E          � � �� n     �  ~h  ��   ��  q
       ���            B  �  �  �         ����  G H          �  �� o     �  �i  `�   ��  q       ���            C  �  �  �         ����  J L          � �� p     �  k  �   ��  q       ���            D  �  �  �         ����  P Q          � �� q       \l  P   ��  q       ���            
E  �  �  �         ����  T U          � �� r     *  �m  �#   ��  q       ���            	F  �  �  �         ����  X Z          � �� s     R  �n  @3   ��  q       ���            G  �  �  �         ����  H I          � �� x     �  lz  |7   ��  r
       ���            B  �  �  �         ����  K M          � �� y       �{  �I   ��  r       ���            C  �  �  �         ����  O P          � %�� z     H  <}  \   ��  r       ���            D  �  �  �         ����  T V          � +�� {     w  �~  Tn   ��  r       ���            E  �  �  �         ����  Y Z          � 1�� |     �  �  ��   ��  r       ���            F  �  �  �         ����  ] _          � 7�� }     �  t�  �   ��  r       ���            G  �  �  �         ����  L M          � 7� �     �  ��  @�   ��  s
       ��8            "L  �  �  �         ����  O Q          � =� �       f�  ��   ��  s       ��8            !M  �  �  �         ����  S U          � C� �     K  �  ��   ��  s       ��8             N  �  �  �         ����  Y [          � I� �     �  r�  <   ��  s       ��8            O  �  �  �         ����  ^ _          � O%� �     �  ��  �   ��  s       ��8            P  �  �  �         ����  b d          � U-� �     �  ~�  �,   ��  s       ��8            Q  �  �  �         ����  Q R          U4� �     m  ڢ  Ɗ	   ��  t
       ��[            .L  �  �  �         ����  U V          [<� �     �  ~�  b�	   ��  t       ��[            -M  �  �  �         ����  Y [          aD� �     �  "�  ��	   ��  t       ��[            ,N  �  �  �         ����  ` a          gL� �     *  Ƨ  ��	   ��  t       ��[            +O  �  �  �         ����  d f          mT� �     i  j�  6�	   ��  t       ��[            *P  �  �  �         ����  i k          $s\�     �  �  �
   ��  t       ��[            )Q  �  �  �         ����  T U          &|b�     �  Z�  ��   ��  u
       ��\            ;V  �  �  �         ����  X Y          ,�j�     �  �  ��   ��  u       ��\            :W  �  �  �         ����  \ ^          2�r�     8  ޼  ��   ��  u       ��\            9X  �  �  �         ����  c d          8�z�     �  ��   �   ��  u       ��\            8Y  �  �  �         ����  h i          >�� �     �  b�      ��  u       ��\            7Z  �  �  �         ����  m o          D��&�       $�  @"   ��  u       ��\            6[  �  �  �         ����  9 :          � � Ul       ?  H:  �      �
       ��l            � .  �  �  8         ����  < =          � � \p       U  8;  �       �       ��l            � /  �  �  8         ����  ? @          � � ct       k  (<  h   ��  �       ��l            � 0  �  �  8         ����  C D          � � jx       �  =  �%   ��  �       ��l            � 1  �  �  8         ����  F H          � � q|       �  >  H.   ��  �       ��l            � 2  �  �  8         ����  J K          � � x�       �  �>  �6   ��  �       ��l            � 3  �  �  8         ����  = >          � � ~{       *  �G  h�   ��  �
       ��m           	 � 8  �  �  9         ����  @ A          � � �       E  �H  ��   ��  �       ��m           	 � 9  �  �  9         ����  C D          � � ��       `  �I  ��   ��  �       ��m           	 � :  �  �  9         ����  H I          � � ��       {  �J  �   ��  �       ��m           	 � ;  �  �  9         ����  K M          � � ��       �  �K  ��   ��  �       ��m           	 � <  �  �  9         ����  O Q          � ��       �  �L  $   ��  �       ��m           	 � =  �  �  9         ����  A B          � ��       �	  �V  ·   ��  �
     	  ��           
 8  �  �           ����  D E          � ��       �	  �W  ��   ��  �     	  ��           
 9  �  �           ����  G I          � ��       �	  �X  ��   ��  �     	  ��           
 :  �  �           ����  L N          � ��       �	  
Z  n�   ��  �     	  ��           
 ;  �  �           ����  P R          � ��       
  6[  R�   ��  �     	  ��           
  <  �  �           ����  T V          � ��       )
  b\  6�   ��  �     	  ��           
 � =  �  �           ����  E F          � !�� n     Z  �f  (�   ��  �
     
  ���            B  �  �  �         ����  H J          � '�� o     �  8h  ��   ��  �     
  ���            C  �  �  �         ����  L M          � -�� p     �  �i  �   ��  �     
  ���            D  �  �  �         ����  Q S          � 3�� q     �  �j  �   ��  �     
  ���            
E  �  �  �         ����  U W          � 9�� r     �  l     ��  �     
  ���            	F  �  �  �         ����  Z [          � ?�� s     "  `m  �    ��  �     
  ���            G  �  �  �         ����  I J          � @�� x     �  �x  ,#   ��  �
       ���            B  �  �  �         ����  M N          � F� y     �  Dz  t5   ��  �       ���            C  �  �  �         ����  P R          � L� z       �{  �G   ��  �       ���            D  �  �  �         ����  V X          R� {     C  }  Z   ��  �       ���            E  �  �  �         ����  Z \          X� |     r  |~  Ll   ��  �       ���            F  �  �  �         ����  _ a          ^%� }     �  �  �~   ��  �       ���            G  �  �  �         ����  L M          ^,� �     �  P�  `�   ��  �
       ��=            "L  �  �  �         ����  O Q          d4� �     �  ֍  ��   ��  �       ��=            !M  �  �  �         ����  S U          j<� �       \�  �   ��  �       ��=             N  �  �  �         ����  Y [          pD� �     J  �  \�   ��  �       ��=            O  �  �  �         ����  ^ _          vL� �     �  h�  �   ��  �       ��=            P  �  �  �         ����  b d          $|T� �     �  �     ��  �       ��=            Q  �  �  �         ����  Q R          ,|[� �     1  J�  Vs	   ��  �
       ��g            .L  �  �  �         ����  U V          2�c� �     p  �  �	   ��  �       ��g            -M  �  �  �         ����  Y [          8�k� �     �  ��  ��	   ��  �       ��g            ,N  �  �  �         ����  ` a          >�s� �     �  6�  *�	   ��  �       ��g            +O  �  �  �         ����  d f          D�{� �     -  ڧ  ��	   ��  �       ��g            *P  �  �  �         ����  i k          J���     l  ~�  b�	   ��  �       ��g            )Q  �  �  �         ����  U V          L���     h  ʷ  �|   ��  �
       ��h            ;V  �  �  �         ����  Y [          R���     �  ��  ��   ��  �       ��h            :W  �  �  �         ����  ^ _          X���     �  N�  �   ��  �       ��h            9X  �  �  �         ����  d f          ^���     @  �   �   ��  �       ��h            8Y  �  �  �         ����  i k          d�� �     �  Ҿ   �   ��  �       ��h            7Z  �  �  �         ����  o p          j��&�     �  ��  @	   ��  �       ��h            6[  �  �  �         ����  9 :          � � ;l         �8  x�      :
       ��            � .  �  �  K         ����  < =          � � Bp       1  �9  �       :       ��            � /  �  �  K         ����  ? @          � � It       G  �:  X   ��  :       ��            � 0  �  �  K         ����  C D          � � Px       ]  �;  �   ��  :       ��            � 1  �  �  K         ����  F H          � � W|       s  x<  8    ��  :       ��            � 2  �  �  K         ����  J K          � � ^�       �  h=  �(   ��  :       ��            � 3  �  �  K         ����  = >          � � d{         F  ȼ   ��  ;
     	  ���           	 � 8  �  �  L         ����  @ A          � � k         "G  T�   ��  ;     	  ���           	 � 9  �  �  L         ����  C D          � � r�       8  0H  ��   ��  ;     	  ���           	 � :  �  �  L         ����  H I          � � y�       S  >I  l�   ��  ;     	  ���           	 � ;  �  �  L         ����  K M          � � ��       n  LJ  ��   ��  ;     	  ���           	 � <  �  �  L         ����  O Q          � � ��       �  ZK  ��   ��  ;     	  ���           	 � =  �  �  L         ����  ? A          � � ��       X	  �T  ��   ��  <
     
  ��!           
 8  �  �           ����  C D          � � ��       y	  "V  v�   ��  <     
  ��!           
 9  �  �           ����  F G          � � ��       �	  NW  Z�   ��  <     
  ��!           
 :  �  �           ����  K L          � � ��       �	  zX  >�   ��  <     
  ��!           
 ;  �  �           ����  O P          � � ��       �	  �Y  "�   ��  <     
  ��!           
  <  �  �           ����  S T          �  ��       �	  �Z  �   ��  <     
  ��!           
 � =  �  �           ����  D E          � �� n     *  ^e  h�   ��  =
       ���            B  �  �  �         ����  G H          � �� o     R  �f  ��   ��  =       ���            C  �  �  �         ����  J L          � �� p     z  �g  X�   ��  =       ���            D  �  �  �         ����  P Q          � �� q     �  <i  ��   ��  =       ���            
E  �  �  �         ����  T U          � �� r     �  �j  H�   ��  =       ���            	F  �  �  �         ����  X Z          � %�� s     �  �k  �   ��  =       ���            G  �  �  �         ����  H I          � &�� x     �  Lw  �   ��  >
       ���            B  �  �  �         ����  K M          � ,�� y     �  �x  $!   ��  >       ���            C  �  �  �         ����  O P          � 2�� z     �  z  l3   ��  >       ���            D  �  �  �         ����  T V          � 8�� {       �{  �E   ��  >       ���            E  �  �  �         ����  Y Z          � >� |     >  �|  �W   ��  >       ���            F  �  �  �         ����  ] _          � D� }     m  T~  Dj   ��  >       ���            G  �  �  �         ����  L M          � D� �     m  ��  ��   ��  ?
       ��B            "L  �  �  �         ����  O Q          � J� �     �  F�  ԫ   ��  ?       ��B            !M  �  �  �         ����  S U          � P"� �     �  ̍  (�   ��  ?       ��B             N  �  �  �         ����  Y [          V*� �       R�  |�   ��  ?       ��B            O  �  �  �         ����  ^ _          \2� �     I  ؐ  ��   ��  ?       ��B            P  �  �  �         ����  b d          b:� �     �  ^�  $   ��  ?       ��B            Q  �  �  �         ����  Q R          bA� �     �  ��  �[	   ��  @
       ��s            .L  �  �           ����  U V          hI� �     4  ^�  �t	   ��  @       ��s            -M  �  �           ����  Y [          nQ� �     s  �  �	   ��  @       ��s            ,N  �  �           ����  ` a          %tY� �     �  ��  ��	   ��  @       ��s            +O  �  �           ����  d f          +za� �     �  J�  V�	   ��  @       ��s            *P  �  �           ����  i k          1�i�     0  �  ��	   ��  @       ��s            )Q  �  �           ����  T U          3�o�     (  :�  �c   ��  A
       ��t            ;V  �  �           ����  X Y          9�w�     p  ��  �   ��  A       ��t            :W  �  �           ����  \ ^          ?��     �  ��  ��   ��  A       ��t            9X  �  �           ����  c d          E���        ��   �   ��  A       ��t            8Y  �  �           ����  h i          K�� �     H  B�   �   ��  A       ��t            7Z  �  �           ����  m o          Q��&�     �  �  @�   ��  A       ��t            6[  �  �           ����  9 :          � � Ml       �  h=  �(      �
     �   �            � .  �  �  ^         ����  < =          � � Tp       �  X>  1       �     �   �            � /  �  �  ^         ����  ? @          � � [t       �  H?  �9   ��  �     �   �            � 0  �  �  ^         ����  C D          � � bx       �  8@  �A   ��  �     �   �            � 1  �  �  ^         ����  F H          � � i|       �  (A  hJ   ��  �     �   �            � 2  �  �  ^         ����  J K          � � p�       �  B  �R   ��  �     �   �            � 3  �  �  ^         ����  = >          � � v{       z  �J  ��   ��  �
     �   �           	 � 8  �  �  _         ����  @ A          � � }       �  �K  4�   ��  �     �   �           	 � 9  �  �  _         ����  C D          � � ��       �  �L  �    ��  �     �   �           	 � :  �  �  _         ����  H I          � � ��       �  �M  L   ��  �     �   �           	 � ;  �  �  _         ����  K M          � � ��       �  �N  �   ��  �     �   �           	 � <  �  �  _         ����  O Q          � � ��         
P  d    ��  �     �   �           	 � =  �  �  _         ����  A B          � � ��       �	  �Y  "�   ��  �
     �   �           
 8  �  �  �         ����  D E          � � ��       �	  �Z  �   ��  �     �   �           
 9  �  �  �         ����  G I          � ��       
  �[  ��   ��  �     �   �           
 :  �  �  �         ����  L N          � ��       ?
  *]  �    ��  �     �   �           
 ;  �  �  �         ����  P R          � ��       `
  V^  �   ��  �     �   �           
  <  �  �  �         ����  T V          � ��       �
  �_  �   ��  �     �   �           
 � =  �  �  �         ����  E F          � �� n     �  j  ��   ��  �
     �   �            B  �  �  �         ����  H J          � �� o     �  Xk      ��  �     �   �            C  �  �  �         ����  L M          � %�� p     
  �l  �   ��  �     �   �            D  �  �  �         ����  Q S          � +�� q     2  �m  '   ��  �     �   �            
E  �  �  �         ����  U W          � 1�� r     Z  6o  �6   ��  �     �   �            	F  �  �  �         ����  Z [          � 7�� s     �  �p   F   ��  �     �   �            G  �  �  �         ����  I J          � 8�� x       �{  �K   ��  �
     �   �            B  �  �  �         ����  M N          � >�� y     M  d}  ^   ��  �     �   �            C  �  �  �         ����  P R          � D� z     |  �~  \p   ��  �     �   �            D  �  �  �         ����  V X          � J� {     �  4�  ��   ��  �     �   �            E  �  �  �         ����  Z \           P� |     �  ��  �   ��  �     �   �            F  �  �  �         ����  _ a          V� }     	  �  4�   ��  �     �   �            G  �  �  �         ����  L M          V$� �       p�   �   ��  �
     �   G            "L  �  �  �         ����  O Q          \,� �     L  ��  t�   ��  �     �   G            !M  �  �  �         ����  S U          b4� �     �  |�  �   ��  �     �   G             N  �  �  �         ����  Y [          h<� �     �  �     ��  �     �   G            O  �  �  �         ����  ^ _          nD� �     �  ��  p-   ��  �     �   G            P  �  �  �         ����  b d          tL� �     (  �  �B   ��  �     �   G            Q  �  �  �         ����  Q R          $tS� �     �  j�  6�	   ��  �
     �               .L  �  �           ����  U V          *z[� �     �  �  Һ	   ��  �     �               -M  �  �           ����  Y [          0�c� �     '  ��  n�	   ��  �     �               ,N  �  �           ����  ` a          6�k� �     f  V�  
�	   ��  �     �               +O  �  �           ����  d f          <�s� �     �  ��  �
   ��  �     �               *P  �  �           ����  i k          B�{�     �  ��  B
   ��  �     �               )Q  �  �           ����  U V          D���     �  �  ��   ��  �
     �   �            ;V  �  �           ����  Y [          J���     0  ��  ��   ��  �     �   �            :W  �  �           ����  ^ _          P���     x  n�  ��   ��  �     �   �            9X  �  �           ����  d f          V���     �  0�      ��  �     �   �            8Y  �  �           ����  i k          \�� �       ��      ��  �     �   �            7Z  �  �           ����  o p          b��&�     P  ��  @;   ��  �     �   �            6[  �  �           ����   9 :          e g       �  (7  h�      E
       ��            � .  �  �  �          ����   < =          i k         8  ��       E       ��            � /  �  �  �          ����   ? @          m o       #  9  H   ��  E       ��            � 0  �  �  �          ����   C D          $q $s       9  �9  �	   ��  E       ��            � 1  �  �  �          ����   F H          *u *w       O  �:  (   ��  E       ��            � 2  �  �  �          ����   J K          0y 0{       e  �;  �   ��  E       ��            � 3  �  �  �          ����   = >          2t 2v       �  �D  (�   ��  F
     	  ��           	 � 8  �  �  �          ����   @ A          8x 8z       �  �E  ��   ��  F     	  ��           	 � 9  �  �  �          ����   C D          >| >~         �F  @�   ��  F     	  ��           	 � :  �  �  �          ����   H I          D� D�       +  �G  ��   ��  F     	  ��           	 � ;  �  �  �          ����   K M          J� J�       F  �H  X�   ��  F     	  ��           	 � <  �  �  �          ����   O Q          P� P�       a  �I  ��   ��  F     	  ��           	 � =  �  �  �          ����   ? A          R� R�       ,	  fS  b�   ��  G
     
  ��           
 8  �  �  �         ����   C D          X� X�       M	  �T  F�   ��  G     
  ��           
 9  �  �  �         ����   F G          ^� ^�       n	  �U  *�   ��  G     
  ��           
 :  �  �  �         ����   K L          d� d�       �	  �V  �   ��  G     
  ��           
 ;  �  �  �         ����   O P          j� j�       �	  X  ��   ��  G     
  ��           
  <  �  �  �         ����   S T          p� p�       �	  BY  ��   ��  G     
  ��           
 � =  �  �  �         ����   D E          {� {� n     �  �c  ��   ��  H
       ���            B  �  �  �         ����   G H          �� �� o     "  e   �   ��  H       ���            C  �  �  �         ����   J L          �� �� p     J  bf  ��   ��  H       ���            D  �  �  �         ����   P Q          �� �� q     r  �g  �   ��  H       ���            
E  �  �  �         ����   T U          �� �� r     �  �h  ��   ��  H       ���            	F  �  �  �         ����   X Z          �� �� s     �  @j   �   ��  H       ���            G  �  �  �         ����   H I          �� �� x     N  �u  ��   ��  I
       ���            B  �  �  �         ����   K M          �� �� y     }  $w  �   ��  I       ���            C  �  �  �         ����   O P          �� �� z     �  �x     ��  I       ���            D  �  �  �         ����   T V          �� �� {     �  �y  d1   ��  I       ���            E  �  �  �         ����   Y Z          �� �� |     
  \{  �C   ��  I       ���            F  �  �  �         ����   ] _          �� �� }     9  �|  �U   ��  I       ���            G  �  �  �         ����   L M          �� �� �     5  0�  ��   ��  J
       ��)            "L  �  �  �         ����   O Q          �� �� �     l  ��  ��   ��  J       ��)            !M  �  �  �         ����   S U          �� �� �     �  <�  H�   ��  J       ��)             N  �  �  �         ����   Y [          �� �� �     �    ��   ��  J       ��)            O  �  �  �         ����   ^ _          �� �� �       H�  ��   ��  J       ��)            P  �  �  �         ����   b d          �� �� �     H  ΐ  D�   ��  J       ��)            Q  �  �  �         ����   Q R          �� �� �     �  *�  vD	   ��  K
       ��9            .L  �  �  �         ����   U V          �� �� �     �  Ο  ]	   ��  K       ��9            -M  �  �  �         ����   Y [          �� �� �     7  r�  �u	   ��  K       ��9            ,N  �  �  �         ����   ` a          � � �     v  �  J�	   ��  K       ��9            +O  �  �  �         ����   d f          � � �     �  ��  �	   ��  K       ��9            *P  �  �  �         ����   i k          � � �     �  ^�  ��	   ��  K       ��9            )Q  �  �  �         ����   T U          !!�     �  ��  �J   ��  L
       ��:            ;V  �  �  �         ����   X Y          ))	�     0  l�  �f   ��  L       ��:            :W  �  �  �         ����   \ ^          11�     x  .�  ��   ��  L       ��:            9X  �  �  �         ����   c d          99�     �  �   �   ��  L       ��:            8Y  �  �  �         ����   h i          AA�       ��   �   ��  L       ��:            7Z  �  �  �         ����   m o          II!�     P  t�  @�   ��  L       ��:            6[  �  �  �         ����  7 9          � e � g       �  45  ��      �
       ��)            � .  �  �  �          ����  : <          i k       �  $6  D�       �       ��)            � /  �  �  �          ����  = ?          	m 	o       �  7  ��   ��  �       ��)            � 0  �  �  �          ����  A C          q s         8  $�   ��  �       ��)            � 1  �  �  �          ����  E F          u w       "  �8  �    ��  �       ��)            � 2  �  �  �          ����  H J          y {       8  �9  	   ��  �       ��)            � 3  �  �  �          ����  ; =          t v       �  �B  ��   ��  �
     	  ��*           	 � 8  �  �  �          ����  > @          #x #z       �  �C  ,�   ��  �     	  ��*           	 � 9  �  �  �          ����  A C          )| )~       �  �D  ��   ��  �     	  ��*           	 � :  �  �  �          ����  F H          /� /�       �  �E  D�   ��  �     	  ��*           	 � ;  �  �  �          ����  J K          5� 5�         �F  ��   ��  �     	  ��*           	 � <  �  �  �          ����  M O          ;� ;�       /  �G  \�   ��  �     	  ��*           	 � =  �  �  �          ����  ? A          =� =�       �  rQ  �   ��  �
     
  ��           
 8  �  �  �         ����  C D          C� C�       	  �R  ʌ   ��  �     
  ��           
 9  �  �  �         ����  F G          I� I�       7	  �S  ��   ��  �     
  ��           
 :  �  �  �         ����  K L          O� O�       X	  �T  ��   ��  �     
  ��           
 ;  �  �  �         ����  O P          U� U�       y	  "V  v�   ��  �     
  ��           
  <  �  �  �         ����  S T          [� [�       �	  NW  Z�   ��  �     
  ��           
 � =  �  �  �         ����  B D          f� f� n     �  �a  8�   ��  �
       ���            B  �  �  �         ����  E G          m� m� o     �  $c  ��   ��  �       ���            C  �  �  �         ����  I J          t� t� p       nd  (�   ��  �       ���            D  �  �  �         ����  N P          {� {� q     6  �e  ��   ��  �       ���            
E  �  �  �         ����  R T          �� �� r     ^  g  �   ��  �       ���            	F  �  �  �         ����  V X          �� �� s     �  Lh  ��   ��  �       ���            G  �  �  �         ����  F H          �� �� x       �s  (�   ��  �
       ���            B  �  �  �         ����  J K          �� �� y     <  0u  p�   ��  �       ���            C  �  �  �         ����  M O          �� �� z     k  �v  �   ��  �       ���            D  �  �  �         ����  S T          �� �� {     �   x      ��  �       ���            E  �  �  �         ����  W Y          �� �� |     �  hy  H*   ��  �       ���            F  �  �  �         ����  [ ]          �� �� }     �  �z  �<   ��  �       ���            G  �  �  �         ����  J L          �� �� �     �  <�  He   ��  �
       ��.            "L  �  �  �         ����  N O          �� �� �     &    �z   ��  �       ��.            !M  �  �  �         ����  R S          �� �� �     ]  H�  ��   ��  �       ��.             N  �  �  �         ����  X Y          �� �� �     �  ΋  D�   ��  �       ��.            O  �  �  �         ����  \ ^          �� �� �     �  T�  ��   ��  �       ��.            P  �  �  �         ����  a b          �� �� �       ڎ  ��   ��  �       ��.            Q  �  �  �         ����  P Q          �� �� �     n  6�  *'	   ��  �
       ��E            .L  �  �  �         ����  T U          �� �� �     �  ڝ  �?	   ��  �       ��E            -M  �  �  �         ����  X Y          �� �� �     �  ~�  bX	   ��  �       ��E            ,N  �  �  �         ����  ^ `          �� �� �     +  "�  �p	   ��  �       ��E            +O  �  �  �         ����  c d          �� �� �     j  Ƣ  ��	   ��  �       ��E            *P  �  �  �         ����  h i          �� �� �     �  j�  6�	   ��  �       ��E            )Q  �  �  �         ����  T U          �     �  ��  `+   ��  �
       ��F            ;V  �  �  �         ����  X Y          	�     �  x�  �G   ��  �       ��F            :W  �  �  �         ����  \ ^          �     (  :�  �c   ��  �       ��F            9X  �  �  �         ����  c d          $$�     p  ��  �   ��  �       ��F            8Y  �  �  �         ����  h i          ,,�     �  ��  ��   ��  �       ��F            7Z  �  �  �         ����  m o          44!�        ��   �   ��  �       ��F            6[  �  �  �         ����  7 9          
e 
g       �  �4  P�      
       ��O            � .  �  �           ����  : <          i k       �  �5  ��              ��O            � /  �  �           ����  = ?          m o       �  �6  0�   ��         ��O            � 0  �  �           ����  A C          q s         �7  ��   ��         ��O            � 1  �  �           ����  E F          "u "w         �8  �   ��         ��O            � 2  �  �           ����  H J          (y ({       /  �9  �   ��         ��O            � 3  �  �           ����  ; =          *t *v       �  ,B  ��   ��  
     	  ��P           	 � 8  �  �           ����  > @          0x 0z       �  :C  D�   ��       	  ��P           	 � 9  �  �           ����  A C          6| 6~       �  HD  Ъ   ��       	  ��P           	 � :  �  �           ����  F H          <� <�       �  VE  \�   ��       	  ��P           	 � ;  �  �           ����  J K          B� B�       
  dF  �   ��       	  ��P           	 � <  �  �           ����  M O          H� H�       %  rG  t�   ��       	  ��P           	 � =  �  �           ����  ? A          J� J�       �  Q  �{   ��  
     
  ��           
 8  �  �  �         ����  C D          P� P�       	  :R  ~�   ��       
  ��           
 9  �  �  �         ����  F G          V� V�       ,	  fS  b�   ��       
  ��           
 :  �  �  �         ����  K L          \� \�       M	  �T  F�   ��       
  ��           
 ;  �  �  �         ����  O P          b� b�       n	  �U  *�   ��       
  ��           
  <  �  �  �         ����  S T          h� h�       �	  �V  �   ��       
  ��           
 � =  �  �  �         ����  B D          s� s� n     �  va  ��   ��  
       ���            B  �  �  �         ����  E G          z� z� o     �  �b   �   ��         ���            C  �  �  �         ����  I J          �� �� p       
d  x�   ��         ���            D  �  �  �         ����  N P          �� �� q     *  Te  �   ��         ���            
E  �  �  �         ����  R T          �� �� r     R  �f  h�   ��         ���            	F  �  �  �         ����  V X          �� �� s     z  �g  ��   ��         ���            G  �  �  �         ����  F H          �� �� x        ds  �   ��  
       ���            B  �  �  �         ����  J K          �� �� y     /  �t  \�   ��         ���            C  �  �  �         ����  M O          �� �� z     ^  4v  �    ��         ���            D  �  �  �         ����  S T          �� �� {     �  �w  �   ��         ���            E  �  �  �         ����  W Y          �� �� |     �  y  4%   ��         ���            F  �  �  �         ����  [ ]          �� �� }     �  lz  |7   ��         ���            G  �  �  �         ����  J L          �� �� �     �  ؆  �_   ��  
       ��4            "L  �  �  �         ����  N O          �� �� �       ^�  $u   ��         ��4            !M  �  �  �         ����  R S          �� �� �     O  �  x�   ��         ��4             N  �  �  �         ����  X Y          �� �� �     �  j�  ̟   ��         ��4            O  �  �  �         ����  \ ^          �� �� �     �  ��   �   ��         ��4            P  �  �  �         ����  a b          �� �� �     �  v�  t�   ��         ��4            Q  �  �  �         ����  P Q          �� �� �     _  қ  N!	   ��  
       ��Q            .L  �  �  �         ����  T U          �� �� �     �  v�  �9	   ��         ��Q            -M  �  �  �         ����  X Y          �� �� �     �  �  �R	   ��         ��Q            ,N  �  �  �         ����  ^ `          �� �� �       ��  "k	   ��         ��Q            +O  �  �  �         ����  c d          � � �     [  b�  ��	   ��         ��Q            *P  �  �  �         ����  h i          � � �     �  �  Z�	   ��         ��Q            )Q  �  �  �         ����  T U          �     �  R�   %   ��   
       ��R            ;V  �  �  �         ����  X Y          !!	�     �  �  @A   ��          ��R            :W  �  �  �         ����  \ ^          ))�       ֵ  `]   ��          ��R            9X  �  �  �         ����  c d          11�     `  ��  �y   ��          ��R            8Y  �  �  �         ����  h i          99�     �  Z�  ��   ��          ��R            7Z  �  �  �         ����  m o          AA!�     �  �  ��   ��          ��R            6[  �  �  �         ����  7 9          � e � g       c  �;  �      
       ��b            � .  �  �  .         ����  : <          � i � k       y  �<  #              ��b            � /  �  �  .         ����  = ?          m o       �  �=  x+   ��         ��b            � 0  �  �  .         ����  A C          
q 
s       �  �>  �3   ��         ��b            � 1  �  �  .         ����  E F          u w       �  �?  X<   ��         ��b            � 2  �  �  .         ����  H J          y {       �  �@  �D   ��         ��b            � 3  �  �  .         ����  ; =          t v       R  4I  �   ��  �
     	  ��c           	 � 8  �  �  /         ����  > @          x z       m  BJ  ��   ��  �     	  ��c           	 � 9  �  �  /         ����  A C          $| $~       �  PK   �   ��  �     	  ��c           	 � :  �  �  /         ����  F H          *� *�       �  ^L  ��   ��  �     	  ��c           	 � ;  �  �  /         ����  J K          0� 0�       �  lM  8   ��  �     	  ��c           	 � <  �  �  /         ����  M O          6� 6�       �  zN  �   ��  �     	  ��c           	 � =  �  �  /         ����  ? A          8� 8�       �	  X  ��   ��  �
     
  ��           
 8  �  �           ����  C D          >� >�       �	  BY  ��   ��  �     
  ��           
 9  �  �           ����  F G          D� D�       �	  nZ  ��   ��  �     
  ��           
 :  �  �           ����  K L          J� J�       
  �[  ��   ��  �     
  ��           
 ;  �  �           ����  O P          P� P�       4
  �\  ��   ��  �     
  ��           
  <  �  �           ����  S T          V� V�       U
  �]  f	   ��  �     
  ��           
 � =  �  �           ����  B D          a� a� n     �  ~h  ��   ��  �
       ���            B  �  �  �         ����  E G          h� h� o     �  �i  `�   ��  �       ���            C  �  �  �         ����  I J          o� o� p     �  k  �   ��  �       ���            D  �  �  �         ����  N P          v� v� q       \l  P   ��  �       ���            
E  �  �  �         ����  R T          }� }� r     *  �m  �#   ��  �       ���            	F  �  �  �         ����  V X          �� �� s     R  �n  @3   ��  �       ���            G  �  �  �         ����  F H          �� �� x     �  lz  |7   ��  �
       ���            B  �  �  �         ����  J K          �� �� y       �{  �I   ��  �       ���            C  �  �  �         ����  M O          �� �� z     H  <}  \   ��  �       ���            D  �  �  �         ����  S T          �� �� {     w  �~  Tn   ��  �       ���            E  �  �  �         ����  W Y          �� �� |     �  �  ��   ��  �       ���            F  �  �  �         ����  [ ]          �� �� }     �  t�  �   ��  �       ���            G  �  �  �         ����  J L          �� �� �     �  ��  @�   ��  �
       ��9            "L  �  �  �         ����  N O          �� �� �       f�  ��   ��  �       ��9            !M  �  �  �         ����  R S          �� �� �     K  �  ��   ��  �       ��9             N  �  �  �         ����  X Y          �� �� �     �  r�  <   ��  �       ��9            O  �  �  �         ����  \ ^          �� �� �     �  ��  �   ��  �       ��9            P  �  �  �         ����  a b          �� �� �     �  ~�  �,   ��  �       ��9            Q  �  �  �         ����  P Q          �� �� �     m  ڢ  Ɗ	   ��  �
       ��]            .L  �  �  �         ����  T U          �� �� �     �  ~�  b�	   ��  �       ��]            -M  �  �  �         ����  X Y          �� �� �     �  "�  ��	   ��  �       ��]            ,N  �  �  �         ����  ^ `          �� �� �     *  Ƨ  ��	   ��  �       ��]            +O  �  �  �         ����  c d          �� �� �     i  j�  6�	   ��  �       ��]            *P  �  �  �         ����  h i          �� �� �     �  �  �
   ��  �       ��]            )Q  �  �  �         ����  T U          �     �  Z�  ��   ��  �
       ��^            ;V  �  �  �         ����  X Y          	�     �  �  ��   ��  �       ��^            :W  �  �  �         ����  \ ^          �     8  ޼  ��   ��  �       ��^            9X  �  �  �         ����  c d          �     �  ��   �   ��  �       ��^            8Y  �  �  �         ����  h i          ''�     �  b�      ��  �       ��^            7Z  �  �  �         ����  m o          //!�       $�  @"   ��  �       ��^            6[  �  �  �         ����  9 :          e g       ?  H:  �      �
       ��u            � .  �  �  A         ����  < =          %i %k       U  8;  �       �       ��u            � /  �  �  A         ����  ? @          +m +o       k  (<  h   ��  �       ��u            � 0  �  �  A         ����  C D          1q 1s       �  =  �%   ��  �       ��u            � 1  �  �  A         ����  F H          7u 7w       �  >  H.   ��  �       ��u            � 2  �  �  A         ����  J K          =y ={       �  �>  �6   ��  �       ��u            � 3  �  �  A         ����  = >          ?t ?v       *  �G  h�   ��  �
       ��v           	 � 8  �  �  B         ����  @ A          Ex Ez       E  �H  ��   ��  �       ��v           	 � 9  �  �  B         ����  C D          K| K~       `  �I  ��   ��  �       ��v           	 � :  �  �  B         ����  H I          Q� Q�       {  �J  �   ��  �       ��v           	 � ;  �  �  B         ����  K M          W� W�       �  �K  ��   ��  �       ��v           	 � <  �  �  B         ����  O Q          ]� ]�       �  �L  $   ��  �       ��v           	 � =  �  �  B         ����  ? A          _� _�       �	  �V  ·   ��  �
     	  ��           
 8  �  �           ����  C D          e� e�       �	  �W  ��   ��  �     	  ��           
 9  �  �           ����  F G          k� k�       �	  �X  ��   ��  �     	  ��           
 :  �  �           ����  K L          q� q�       �	  
Z  n�   ��  �     	  ��           
 ;  �  �           ����  O P          w� w�       
  6[  R�   ��  �     	  ��           
  <  �  �           ����  S T          }� }�       )
  b\  6�   ��  �     	  ��           
 � =  �  �           ����  D E          �� �� n     Z  �f  (�   ��  �
     
  ���            B  �  �  �         ����  G H          �� �� o     �  8h  ��   ��  �     
  ���            C  �  �  �         ����  J L          �� �� p     �  �i  �   ��  �     
  ���            D  �  �  �         ����  P Q          �� �� q     �  �j  �   ��  �     
  ���            
E  �  �  �         ����  T U          �� �� r     �  l     ��  �     
  ���            	F  �  �  �         ����  X Z          �� �� s     "  `m  �    ��  �     
  ���            G  �  �  �         ����  H I          �� �� x     �  �x  ,#   ��  �
       ���            B  �  �  �         ����  K M          �� �� y     �  Dz  t5   ��  �       ���            C  �  �  �         ����  O P          �� �� z       �{  �G   ��  �       ���            D  �  �  �         ����  T V          �� �� {     C  }  Z   ��  �       ���            E  �  �  �         ����  Y Z          �� �� |     r  |~  Ll   ��  �       ���            F  �  �  �         ����  ] _          �� �� }     �  �  �~   ��  �       ���            G  �  �  �         ����  L M          �� �� �     �  P�  `�   ��  �
       ��>            "L  �  �  �         ����  O Q          �� �� �     �  ֍  ��   ��  �       ��>            !M  �  �  �         ����  S U          �� �� �       \�  �   ��  �       ��>             N  �  �  �         ����  Y [          �� �� �     J  �  \�   ��  �       ��>            O  �  �  �         ����  ^ _          �� �� �     �  h�  �   ��  �       ��>            P  �  �  �         ����  b d          �� �� �     �  �     ��  �       ��>            Q  �  �  �         ����  Q R          �� �� �     1  J�  Vs	   ��  �
       ��i            .L  �  �  �         ����  U V          � � �     p  �  �	   ��  �       ��i            -M  �  �  �         ����  Y [          � � �     �  ��  ��	   ��  �       ��i            ,N  �  �  �         ����  ` a          � � �     �  6�  *�	   ��  �       ��i            +O  �  �  �         ����  d f          � � �     -  ڧ  ��	   ��  �       ��i            *P  �  �  �         ����  i k          !� !� �     l  ~�  b�	   ��  �       ��i            )Q  �  �  �         ����  T U          ..�     h  ʷ  �|   ��  �
       ��j            ;V  �  �  �         ����  X Y          66	�     �  ��  ��   ��  �       ��j            :W  �  �  �         ����  \ ^          >>�     �  N�  �   ��  �       ��j            9X  �  �  �         ����  c d          FF�     @  �   �   ��  �       ��j            8Y  �  �  �         ����  h i          NN�     �  Ҿ   �   ��  �       ��j            7Z  �  �  �         ����  m o          VV!�     �  ��  @	   ��  �       ��j            6[  �  �  �         ����  7 9          e g         �8  x�      K
       ���            � .  �  �  T         ����  : <          i k       1  �9  �       K       ���            � /  �  �  T         ����  = ?          m o       G  �:  X   ��  K       ���            � 0  �  �  T         ����  A C          q s       ]  �;  �   ��  K       ���            � 1  �  �  T         ����  E F          u w       s  x<  8    ��  K       ���            � 2  �  �  T         ����  H J          #y #{       �  h=  �(   ��  K       ���            � 3  �  �  T         ����  ; =          %t %v         F  ȼ   ��  L
     	  ���           	 � 8  �  �  U         ����  > @          +x +z         "G  T�   ��  L     	  ���           	 � 9  �  �  U         ����  A C          1| 1~       8  0H  ��   ��  L     	  ���           	 � :  �  �  U         ����  F H          7� 7�       S  >I  l�   ��  L     	  ���           	 � ;  �  �  U         ����  J K          =� =�       n  LJ  ��   ��  L     	  ���           	 � <  �  �  U         ����  M O          C� C�       �  ZK  ��   ��  L     	  ���           	 � =  �  �  U         ����  ? A          E� E�       X	  �T  ��   ��  M
     
  ��#           
 8  �  �           ����  C D          K� K�       y	  "V  v�   ��  M     
  ��#           
 9  �  �           ����  F G          Q� Q�       �	  NW  Z�   ��  M     
  ��#           
 :  �  �           ����  K L          W� W�       �	  zX  >�   ��  M     
  ��#           
 ;  �  �           ����  O P          ]� ]�       �	  �Y  "�   ��  M     
  ��#           
  <  �  �           ����  S T          c� c�       �	  �Z  �   ��  M     
  ��#           
 � =  �  �           ����  B D          n� n� n     *  ^e  h�   ��  N
       ���            B  �  �  �         ����  E G          u� u� o     R  �f  ��   ��  N       ���            C  �  �  �         ����  I J          |� |� p     z  �g  X�   ��  N       ���            D  �  �  �         ����  N P          �� �� q     �  <i  ��   ��  N       ���            
E  �  �  �         ����  R T          �� �� r     �  �j  H�   ��  N       ���            	F  �  �  �         ����  V X          �� �� s     �  �k  �   ��  N       ���            G  �  �  �         ����  F H          �� �� x     �  Lw  �   ��  O
       ���            B  �  �  �         ����  J K          �� �� y     �  �x  $!   ��  O       ���            C  �  �  �         ����  M O          �� �� z     �  z  l3   ��  O       ���            D  �  �  �         ����  S T          �� �� {       �{  �E   ��  O       ���            E  �  �  �         ����  W Y          �� �� |     >  �|  �W   ��  O       ���            F  �  �  �         ����  [ ]          �� �� }     m  T~  Dj   ��  O       ���            G  �  �  �         ����  J L          �� �� �     m  ��  ��   ��  P
       ��C            "L  �  �  �         ����  N O          �� �� �     �  F�  ԫ   ��  P       ��C            !M  �  �  �         ����  R S          �� �� �     �  ̍  (�   ��  P       ��C             N  �  �  �         ����  X Y          �� �� �       R�  |�   ��  P       ��C            O  �  �  �         ����  \ ^          �� �� �     I  ؐ  ��   ��  P       ��C            P  �  �  �         ����  a b          �� �� �     �  ^�  $   ��  P       ��C            Q  �  �  �         ����  P Q          �� �� �     �  ��  �[	   ��  Q
       ��u            .L  �  �           ����  T U          �� �� �     4  ^�  �t	   ��  Q       ��u            -M  �  �           ����  X Y          �� �� �     s  �  �	   ��  Q       ��u            ,N  �  �           ����  ^ `          �� �� �     �  ��  ��	   ��  Q       ��u            +O  �  �           ����  c d           �  � �     �  J�  V�	   ��  Q       ��u            *P  �  �           ����  h i          � � �     0  �  ��	   ��  Q       ��u            )Q  �  �           ����  Q R          �     (  :�  �c   ��  R
       ��v            ;V  �  �  	         ����  U V          	�     p  ��  �   ��  R       ��v            :W  �  �  	         ����  Y [          $$�     �  ��  ��   ��  R       ��v            9X  �  �  	         ����  ` a          ,,�        ��   �   ��  R       ��v            8Y  �  �  	         ����  d f          44�     H  B�   �   ��  R       ��v            7Z  �  �  	         ����  i k          <<!�     �  �  @�   ��  R       ��v            6[  �  �  	         ����  9 :          e g       �  h=  �(      �
     �   �            � .  �  �  g         ����  < =          i k       �  X>  1       �     �   �            � /  �  �  g         ����  ? @          #m #o       �  H?  �9   ��  �     �   �            � 0  �  �  g         ����  C D          )q )s       �  8@  �A   ��  �     �   �            � 1  �  �  g         ����  F H          /u /w       �  (A  hJ   ��  �     �   �            � 2  �  �  g         ����  J K          5y 5{       �  B  �R   ��  �     �   �            � 3  �  �  g         ����  = >          7t 7v       z  �J  ��   ��  �
     �   �           	 � 8  �  �  h         ����  @ A          =x =z       �  �K  4�   ��  �     �   �           	 � 9  �  �  h         ����  C D          C| C~       �  �L  �    ��  �     �   �           	 � :  �  �  h         ����  H I          I� I�       �  �M  L   ��  �     �   �           	 � ;  �  �  h         ����  K M          O� O�       �  �N  �   ��  �     �   �           	 � <  �  �  h         ����  O Q          U� U�         
P  d    ��  �     �   �           	 � =  �  �  h         ����  ? A          W� W�       �	  �Y  "�   ��  �
     �   �           
 8  �  �  �         ����  C D          ]� ]�       �	  �Z  �   ��  �     �   �           
 9  �  �  �         ����  F G          c� c�       
  �[  ��   ��  �     �   �           
 :  �  �  �         ����  K L          i� i�       ?
  *]  �    ��  �     �   �           
 ;  �  �  �         ����  O P          o� o�       `
  V^  �   ��  �     �   �           
  <  �  �  �         ����  S T          u� u�       �
  �_  �   ��  �     �   �           
 � =  �  �  �         ����  D E          �� �� n     �  j  ��   ��  �
     �   �            B  �  �  �         ����  G H          �� �� o     �  Xk      ��  �     �   �            C  �  �  �         ����  J L          �� �� p     
  �l  �   ��  �     �   �            D  �  �  �         ����  P Q          �� �� q     2  �m  '   ��  �     �   �            
E  �  �  �         ����  T U          �� �� r     Z  6o  �6   ��  �     �   �            	F  �  �  �         ����  X Z          �� �� s     �  �p   F   ��  �     �   �            G  �  �  �         ����  H I          �� �� x       �{  �K   ��  �
     �   �            B  �  �  �         ����  K M          �� �� y     M  d}  ^   ��  �     �   �            C  �  �  �         ����  O P          �� �� z     |  �~  \p   ��  �     �   �            D  �  �  �         ����  T V          �� �� {     �  4�  ��   ��  �     �   �            E  �  �  �         ����  Y Z          �� �� |     �  ��  �   ��  �     �   �            F  �  �  �         ����  ] _          �� �� }     	  �  4�   ��  �     �   �            G  �  �  �         ����  L M          �� �� �       p�   �   ��  �
     �   H            "L  �  �  �         ����  O Q          �� �� �     L  ��  t�   ��  �     �   H            !M  �  �  �         ����  S U          �� �� �     �  |�  �   ��  �     �   H             N  �  �  �         ����  Y [          �� �� �     �  �     ��  �     �   H            O  �  �  �         ����  ^ _          �� �� �     �  ��  p-   ��  �     �   H            P  �  �  �         ����  b d          �� �� �     (  �  �B   ��  �     �   H            Q  �  �  �         ����  Q R          �� �� �     �  j�  6�	   ��  �
     �   �            .L  �  �           ����  U V          �� �� �     �  �  Һ	   ��  �     �   �            -M  �  �           ����  Y [          � � �     '  ��  n�	   ��  �     �   �            ,N  �  �           ����  ` a          � � �     f  V�  
�	   ��  �     �   �            +O  �  �           ����  d f          � � �     �  ��  �
   ��  �     �   �            *P  �  �           ����  i k          � � �     �  ��  B
   ��  �     �   �            )Q  �  �           ����  T U          &&�     �  �  ��   ��  �
     �   �            ;V  �  �           ����  X Y          ..	�     0  ��  ��   ��  �     �   �            :W  �  �           ����  \ ^          66�     x  n�  ��   ��  �     �   �            9X  �  �           ����  c d          >>�     �  0�      ��  �     �   �            8Y  �  �           ����  h i          FF�       ��      ��  �     �   �            7Z  �  �           ����  m o          NN!�     P  ��  @;   ��  �     �   �            6[  �  �           ����   1 2          { � Jm       �  (7  h�      Y
       ��(            � .  �  �           ����   3 4           � Qq         8  ��       Y       ��(            � /  �  �           ����   6 7          � � Xu       #  9  H   ��  Y       ��(            � 0  �  �           ����   9 ;          � � _y       9  �9  �	   ��  Y       ��(            � 1  �  �           ����   < >          � � f}       O  �:  (   ��  Y       ��(            � 2  �  �           ����   ? A          � � m�       e  �;  �   ��  Y       ��(            � 3  �  �           ����   3 5          � � s|       �  �D  (�   ��  Z
     	  ��)           	 � 8  �  �           ����   6 7          � � z�       �  �E  ��   ��  Z     	  ��)           	 � 9  �  �           ����   9 :          � � ��         �F  @�   ��  Z     	  ��)           	 � :  �  �           ����   = >          � � ��       +  �G  ��   ��  Z     	  ��)           	 � ;  �  �           ����   @ A          � � ��       F  �H  X�   ��  Z     	  ��)           	 � <  �  �           ����   C D          � � ��       a  �I  ��   ��  Z     	  ��)           	 � =  �  �           ����   6 7          � � ��       ,	  fS  b�   ��  [
     
  ��*           
 8  �  �           ����   9 :          � � ��       M	  �T  F�   ��  [     
  ��*           
 9  �  �           ����   < =          � � ��       n	  �U  *�   ��  [     
  ��*           
 :  �  �           ����   @ A          � � ��       �	  �V  �   ��  [     
  ��*           
 ;  �  �           ����   C E          � � ��       �	  X  ��   ��  [     
  ��*           
  <  �  �           ����   F H          � ��       �	  BY  ��   ��  [     
  ��*           
 � =  �  �           ����   : ;          � 	�� n     �  �c  ��   ��  \
       ���            B  �  �  �         ����   = >          � �� o     "  e   �   ��  \       ���            C  �  �  �         ����   @ A          � �� p     J  bf  ��   ��  \       ���            D  �  �  �         ����   D F          � �� q     r  �g  �   ��  \       ���            
E  �  �  �         ����   H J          � !�� r     �  �h  ��   ��  \       ���            	F  �  �  �         ����   K M          � '�� s     �  @j   �   ��  \       ���            G  �  �  �         ����   = >          � (�� x     N  �u  ��   ��  ]
       ���            B  �  �  �         ����   @ A          � .�� y     }  $w  �   ��  ]       ���            C  �  �  �         ����   C D          � 4� z     �  �x     ��  ]       ���            D  �  �  �         ����   H I          � :
� {     �  �y  d1   ��  ]       ���            E  �  �  �         ����   K M          � @� |     
  \{  �C   ��  ]       ���            F  �  �  �         ����   O Q          � F� }     9  �|  �U   ��  ]       ���            G  �  �  �         ����   ? A          � F!� �     5  0�  ��   ��  ^
       ��*            "L  �  �  �         ����   C D          � L)� �     l  ��  ��   ��  ^       ��*            !M  �  �  �         ����   F G          � R1� �     �  <�  H�   ��  ^       ��*             N  �  �  �         ����   K L          � X9� �     �    ��   ��  ^       ��*            O  �  �  �         ����   O P          � ^A� �       H�  ��   ��  ^       ��*            P  �  �  �         ����   S T          dI� �     H  ΐ  D�   ��  ^       ��*            Q  �  �  �         ����   D E          dP� �     �  *�  vD	   ��  _
       ��;            .L  �  �  �         ����   G H          jX� �     �  Ο  ]	   ��  _       ��;            -M  �  �  �         ����   J L          p`� �     7  r�  �u	   ��  _       ��;            ,N  �  �  �         ����   P Q          vh� �     v  �  J�	   ��  _       ��;            +O  �  �  �         ����   T U          #|p� �     �  ��  �	   ��  _       ��;            *P  �  �  �         ����   X Z          )�x�     �  ^�  ��	   ��  _       ��;            )Q  �  �  �         ����   F H          +�~	�     �  ��  �J   ��  `
       ��<            ;V  �  �  �         ����   J K          1���     0  l�  �f   ��  `       ��<            :W  �  �  �         ����   M O          7���     x  .�  ��   ��  `       ��<            9X  �  �  �         ����   S T          =���     �  �   �   ��  `       ��<            8Y  �  �  �         ����   W Y          C��!�       ��   �   ��  `       ��<            7Z  �  �  �         ����   [ ]          I��'�     P  t�  @�   ��  `       ��<            6[  �  �  �         ����  1 2          r � Ad       �  45  ��      �
       ��-            � .  �  �           ����  3 4          v � Hh       �  $6  D�       �       ��-            � /  �  �           ����  6 7          z � Ol       �  7  ��   ��  �       ��-            � 0  �  �           ����  9 ;          ~ � Vp         8  $�   ��  �       ��-            � 1  �  �           ����  < >          � � ]t       "  �8  �    ��  �       ��-            � 2  �  �           ����  ? A          � � dx       8  �9  	   ��  �       ��-            � 3  �  �           ����  3 5          � � js       �  �B  ��   ��  �
     	  ��.           	 � 8  �  �           ����  6 7          � � qw       �  �C  ,�   ��  �     	  ��.           	 � 9  �  �           ����  9 :          � � x{       �  �D  ��   ��  �     	  ��.           	 � :  �  �           ����  = >          � �        �  �E  D�   ��  �     	  ��.           	 � ;  �  �           ����  @ A          � � ��         �F  ��   ��  �     	  ��.           	 � <  �  �           ����  C D          � � ��       /  �G  \�   ��  �     	  ��.           	 � =  �  �           ����  6 7          � � ��       �  rQ  �   ��  �
     
  ��/           
 8  �  �           ����  9 :          � � ��       	  �R  ʌ   ��  �     
  ��/           
 9  �  �           ����  < =          � � ��       7	  �S  ��   ��  �     
  ��/           
 :  �  �           ����  @ A          � � ��       X	  �T  ��   ��  �     
  ��/           
 ;  �  �           ����  C E          � � ��       y	  "V  v�   ��  �     
  ��/           
  <  �  �           ����  F H          � � ��       �	  NW  Z�   ��  �     
  ��/           
 � =  �  �           ����  9 :          �  �� n     �  �a  8�   ��  �
       ���            B  �  �  �         ����  < =          � �� o     �  $c  ��   ��  �       ���            C  �  �  �         ����  ? @          � �� p       nd  (�   ��  �       ���            D  �  �  �         ����  C D          � �� q     6  �e  ��   ��  �       ���            
E  �  �  �         ����  F H          � �� r     ^  g  �   ��  �       ���            	F  �  �  �         ����  J K          � �� s     �  Lh  ��   ��  �       ���            G  �  �  �         ����  ; =          � �� x       �s  (�   ��  �
       ���            B  �  �  �         ����  > @          � %�� y     <  0u  p�   ��  �       ���            C  �  �  �         ����  A C          � +�� z     k  �v  �   ��  �       ���            D  �  �  �         ����  F H          � 1� {     �   x      ��  �       ���            E  �  �  �         ����  J K          � 7	� |     �  hy  H*   ��  �       ���            F  �  �  �         ����  M O          � =� }     �  �z  �<   ��  �       ���            G  �  �  �         ����  > ?          � =� �     �  <�  He   ��  �
       ��/            "L  �  �  �         ����  A C          � C � �     &    �z   ��  �       ��/            !M  �  �  �         ����  D F          � I(� �     ]  H�  ��   ��  �       ��/             N  �  �  �         ����  I K          � O0� �     �  ΋  D�   ��  �       ��/            O  �  �  �         ����  M O          � U8� �     �  T�  ��   ��  �       ��/            P  �  �  �         ����  Q S          � [@� �       ڎ  ��   ��  �       ��/            Q  �  �  �         ����  B D          [G� �     n  6�  *'	   ��  �
       ��G            .L  �  �  �         ����  E G          aO� �     �  ڝ  �?	   ��  �       ��G            -M  �  �  �         ����  I J          gW� �     �  ~�  bX	   ��  �       ��G            ,N  �  �  �         ����  N P          m_� �     +  "�  �p	   ��  �       ��G            +O  �  �  �         ����  R T          sg� �     j  Ƣ  ��	   ��  �       ��G            *P  �  �  �         ����  V X           yo� �     �  j�  6�	   ��  �       ��G            )Q  �  �  �         ����  E F          "�u �     �  ��  `+   ��  �
       ��H            ;V  �  �  �         ����  H J          (�}�     �  x�  �G   ��  �       ��H            :W  �  �  �         ����  L M          .���     (  :�  �c   ��  �       ��H            9X  �  �  �         ����  Q S          4���     p  ��  �   ��  �       ��H            8Y  �  �  �         ����  U W          :���     �  ��  ��   ��  �       ��H            7Z  �  �  �         ����  Z [          @���        ��   �   ��  �       ��H            6[  �  �  �         ����  1 2          � � Dm       �  �4  P�      *
       ��2            � .  �  �           ����  3 4          � � Kq       �  �5  ��       *       ��2            � /  �  �           ����  6 7          � � Ru       �  �6  0�   ��  *       ��2            � 0  �  �           ����  9 ;          � � Yy         �7  ��   ��  *       ��2            � 1  �  �           ����  < >          � � `}         �8  �   ��  *       ��2            � 2  �  �           ����  ? A          � � g�       /  �9  �   ��  *       ��2            � 3  �  �           ����  3 5          � � m|       �  ,B  ��   ��  +
     	  ��3           	 � 8  �  �           ����  6 7          � � t�       �  :C  D�   ��  +     	  ��3           	 � 9  �  �           ����  9 :          � � {�       �  HD  Ъ   ��  +     	  ��3           	 � :  �  �           ����  = >          � � ��       �  VE  \�   ��  +     	  ��3           	 � ;  �  �           ����  @ A          � � ��       
  dF  �   ��  +     	  ��3           	 � <  �  �           ����  C D          � � ��       %  rG  t�   ��  +     	  ��3           	 � =  �  �           ����  6 7          � � ��       �  Q  �{   ��  ,
     
  ��4           
 8  �  �           ����  9 :          � � ��       	  :R  ~�   ��  ,     
  ��4           
 9  �  �           ����  < =          � � ��       ,	  fS  b�   ��  ,     
  ��4           
 :  �  �           ����  @ A          � � ��       M	  �T  F�   ��  ,     
  ��4           
 ;  �  �           ����  C E          � � ��       n	  �U  *�   ��  ,     
  ��4           
  <  �  �           ����  F H          � ��       �	  �V  �   ��  ,     
  ��4           
 � =  �  �           ����  9 :          � �� n     �  va  ��   ��  -
       ���            B  �  �  �         ����  < =          � �� o     �  �b   �   ��  -       ���            C  �  �  �         ����  ? @          � �� p       
d  x�   ��  -       ���            D  �  �  �         ����  C D          � �� q     *  Te  �   ��  -       ���            
E  �  �  �         ����  F H          � #�� r     R  �f  h�   ��  -       ���            	F  �  �  �         ����  J K          � )�� s     z  �g  ��   ��  -       ���            G  �  �  �         ����  ; =          � *�� x        ds  �   ��  .
       ���            B  �  �  �         ����  > @          � 0�� y     /  �t  \�   ��  .       ���            C  �  �  �         ����  A C          � 6�� z     ^  4v  �    ��  .       ���            D  �  �  �         ����  F H          � <� {     �  �w  �   ��  .       ���            E  �  �  �         ����  J K          � B� |     �  y  4%   ��  .       ���            F  �  �  �         ����  M O          � H� }     �  lz  |7   ��  .       ���            G  �  �  �         ����  > ?          � H� �     �  ؆  �_   ��  /
       ��5            "L  �  �  �         ����  A C          � N#� �       ^�  $u   ��  /       ��5            !M  �  �  �         ����  D F          � T+� �     O  �  x�   ��  /       ��5             N  �  �  �         ����  I K          Z3� �     �  j�  ̟   ��  /       ��5            O  �  �  �         ����  M O          `;� �     �  ��   �   ��  /       ��5            P  �  �  �         ����  Q S          fC� �     �  v�  t�   ��  /       ��5            Q  �  �  �         ����  B D          fJ� �     _  қ  N!	   ��  0
       ��S            .L  �  �  �         ����  E G          lR� �     �  v�  �9	   ��  0       ��S            -M  �  �  �         ����  I J           rZ� �     �  �  �R	   ��  0       ��S            ,N  �  �  �         ����  N P          &xb� �       ��  "k	   ��  0       ��S            +O  �  �  �         ����  R T          ,~j� �     [  b�  ��	   ��  0       ��S            *P  �  �  �         ����  V X          2�r�     �  �  Z�	   ��  0       ��S            )Q  �  �  �         ����  E F          4�x	�     �  R�   %   ��  1
       ��T            ;V  �  �  �         ����  H J          :���     �  �  @A   ��  1       ��T            :W  �  �  �         ����  L M          @���       ֵ  `]   ��  1       ��T            9X  �  �  �         ����  Q S          F���     `  ��  �y   ��  1       ��T            8Y  �  �  �         ����  U W          L��!�     �  Z�  ��   ��  1       ��T            7Z  �  �  �         ����  Z [          R��'�     �  �  ��   ��  1       ��T            6[  �  �  �         ����  1 2          o � >a       c  �;  �      �
       ��7            � .  �  �  !         ����  3 4          s � Ee       y  �<  #       �       ��7            � /  �  �  !         ����  6 7          w � Li       �  �=  x+   ��  �       ��7            � 0  �  �  !         ����  9 ;          { � Sm       �  �>  �3   ��  �       ��7            � 1  �  �  !         ����  < >           � Zq       �  �?  X<   ��  �       ��7            � 2  �  �  !         ����  ? A          � � au       �  �@  �D   ��  �       ��7            � 3  �  �  !         ����  3 5          ~ � gp       R  4I  �   ��  �
     	  ��8           	 � 8  �  �  "         ����  6 7          � � nt       m  BJ  ��   ��  �     	  ��8           	 � 9  �  �  "         ����  9 :          � � ux       �  PK   �   ��  �     	  ��8           	 � :  �  �  "         ����  = >          � � ||       �  ^L  ��   ��  �     	  ��8           	 � ;  �  �  "         ����  @ A          � � ��       �  lM  8   ��  �     	  ��8           	 � <  �  �  "         ����  C D          � � ��       �  zN  �   ��  �     	  ��8           	 � =  �  �  "         ����  6 7          � � �       �	  X  ��   ��  �
     
  ��9           
 8  �  �  #         ����  9 :          � � ��       �	  BY  ��   ��  �     
  ��9           
 9  �  �  #         ����  < =          � � ��       �	  nZ  ��   ��  �     
  ��9           
 :  �  �  #         ����  @ A          � � ��       
  �[  ��   ��  �     
  ��9           
 ;  �  �  #         ����  C E          � � ��       4
  �\  ��   ��  �     
  ��9           
  <  �  �  #         ����  F H          � � ��       U
  �]  f	   ��  �     
  ��9           
 � =  �  �  #         ����  9 :          � � �� n     �  ~h  ��   ��  �
       ���            B  �  �  �         ����  < =          � �� o     �  �i  `�   ��  �       ���            C  �  �  �         ����  ? @          � 	�� p     �  k  �   ��  �       ���            D  �  �  �         ����  C D          � �� q       \l  P   ��  �       ���            
E  �  �  �         ����  F H          � �� r     *  �m  �#   ��  �       ���            	F  �  �  �         ����  J K          � �� s     R  �n  @3   ��  �       ���            G  �  �  �         ����  ; =          � �� x     �  lz  |7   ��  �
       ���            B  �  �  �         ����  > @          � "�� y       �{  �I   ��  �       ���            C  �  �  �         ����  A C          � (�� z     H  <}  \   ��  �       ���            D  �  �  �         ����  F H          � .�� {     w  �~  Tn   ��  �       ���            E  �  �  �         ����  J K          � 4� |     �  �  ��   ��  �       ���            F  �  �  �         ����  M O          � :� }     �  t�  �   ��  �       ���            G  �  �  �         ����  > ?          � :� �     �  ��  @�   ��  �
       ��:            "L  �  �  �         ����  A C          � @� �       f�  ��   ��  �       ��:            !M  �  �  �         ����  D F          � F%� �     K  �  ��   ��  �       ��:             N  �  �  �         ����  I K          � L-� �     �  r�  <   ��  �       ��:            O  �  �  �         ����  M O          � R5� �     �  ��  �   ��  �       ��:            P  �  �  �         ����  Q S          � X=� �     �  ~�  �,   ��  �       ��:            Q  �  �  �         ����  B D          � XD� �     m  ڢ  Ɗ	   ��  �
       ��_            .L  �  �  �         ����  E G          ^L� �     �  ~�  b�	   ��  �       ��_            -M  �  �  �         ����  I J          dT� �     �  "�  ��	   ��  �       ��_            ,N  �  �  �         ����  N P          j\� �     *  Ƨ  ��	   ��  �       ��_            +O  �  �  �         ����  R T          pd� �     i  j�  6�	   ��  �       ��_            *P  �  �  �         ����  V X          vl� �     �  �  �
   ��  �       ��_            )Q  �  �  �         ����  E F          r� �     �  Z�  ��   ��  �
       ��`            ;V  �  �  �         ����  H J          %�z�     �  �  ��   ��  �       ��`            :W  �  �  �         ����  L M          +��	�     8  ޼  ��   ��  �       ��`            9X  �  �  �         ����  Q S          1���     �  ��   �   ��  �       ��`            8Y  �  �  �         ����  U W          7���     �  b�      ��  �       ��`            7Z  �  �  �         ����  Z [          =���       $�  @"   ��  �       ��`            6[  �  �  �         ����  1 2          � � Y|       ?  H:  �      �
       ��<            � .  �  �  &         ����  3 4          � � `�       U  8;  �       �       ��<            � /  �  �  &         ����  6 7          � � g�       k  (<  h   ��  �       ��<            � 0  �  �  &         ����  9 ;          � � n�       �  =  �%   ��  �       ��<            � 1  �  �  &         ����  < >          � � u�       �  >  H.   ��  �       ��<            � 2  �  �  &         ����  ? A          � � |�       �  �>  �6   ��  �       ��<            � 3  �  �  &         ����  3 5          � � ��       *  �G  h�   ��  �
       ��=           	 � 8  �  �  '         ����  6 7          � � ��       E  �H  ��   ��  �       ��=           	 � 9  �  �  '         ����  9 :          � � ��       `  �I  ��   ��  �       ��=           	 � :  �  �  '         ����  = >          � � ��       {  �J  �   ��  �       ��=           	 � ;  �  �  '         ����  @ A          � � ��       �  �K  ��   ��  �       ��=           	 � <  �  �  '         ����  C D          � � ��       �  �L  $   ��  �       ��=           	 � =  �  �  '         ����  6 7          � � ��       �	  �V  ·   ��  �
     	  ��>           
 8  �  �  (         ����  9 :          � � ��       �	  �W  ��   ��  �     	  ��>           
 9  �  �  (         ����  < =          � ��       �	  �X  ��   ��  �     	  ��>           
 :  �  �  (         ����  @ A          � ��       �	  
Z  n�   ��  �     	  ��>           
 ;  �  �  (         ����  C E          � ��       
  6[  R�   ��  �     	  ��>           
  <  �  �  (         ����  F H          � ��       )
  b\  6�   ��  �     	  ��>           
 � =  �  �  (         ����  : ;          � �� n     Z  �f  (�   ��  �
     
  ���            B  �  �  �         ����  = >          � �� o     �  8h  ��   ��  �     
  ���            C  �  �  �         ����  @ A          � $�� p     �  �i  �   ��  �     
  ���            D  �  �  �         ����  D F          � *�� q     �  �j  �   ��  �     
  ���            
E  �  �  �         ����  H J          � 0�� r     �  l     ��  �     
  ���            	F  �  �  �         ����  K M          � 6�� s     "  `m  �    ��  �     
  ���            G  �  �  �         ����  = >          � 7� x     �  �x  ,#   ��  �
       ���            B  �  �  �         ����  @ A          � =	� y     �  Dz  t5   ��  �       ���            C  �  �  �         ����  C D          � C� z       �{  �G   ��  �       ���            D  �  �  �         ����  H I          � I� {     C  }  Z   ��  �       ���            E  �  �  �         ����  K M          � O!� |     r  |~  Ll   ��  �       ���            F  �  �  �         ����  O Q          � U)� }     �  �  �~   ��  �       ���            G  �  �  �         ����  ? A          � U0� �     �  P�  `�   ��  �
       ��?            "L  �  �  �         ����  C D          � [8� �     �  ֍  ��   ��  �       ��?            !M  �  �  �         ����  F G          a@� �       \�  �   ��  �       ��?             N  �  �  �         ����  K L          gH� �     J  �  \�   ��  �       ��?            O  �  �  �         ����  O P          mP� �     �  h�  �   ��  �       ��?            P  �  �  �         ����  S T          sX� �     �  �     ��  �       ��?            Q  �  �  �         ����  D E          s_� �     1  J�  Vs	   ��  �
       ��k            .L  �  �  �         ����  G H           yg� �     p  �  �	   ��  �       ��k            -M  �  �  �         ����  J L          &o�     �  ��  ��	   ��  �       ��k            ,N  �  �  �         ����  P Q          ,�w�     �  6�  *�	   ��  �       ��k            +O  �  �  �         ����  T U          2��     -  ڧ  ��	   ��  �       ��k            *P  �  �  �         ����  X Z          8���     l  ~�  b�	   ��  �       ��k            )Q  �  �  �         ����  F H          :���     h  ʷ  �|   ��  �
       ��l            ;V  �  �  �         ����  J K          @���     �  ��  ��   ��  �       ��l            :W  �  �  �         ����  M O          F��$�     �  N�  �   ��  �       ��l            9X  �  �  �         ����  S T          L��*�     @  �   �   ��  �       ��l            8Y  �  �  �         ����  W Y          R��0�     �  Ҿ   �   ��  �       ��l            7Z  �  �  �         ����  [ ]          X��6�     �  ��  @	   ��  �       ��l            6[  �  �  �         ����  1 2          � � Ps         �8  x�      \
       ��A            � .  �  �  +         ����  3 4          � � Ww       1  �9  �       \       ��A            � /  �  �  +         ����  6 7          � � ^{       G  �:  X   ��  \       ��A            � 0  �  �  +         ����  9 ;          � � e       ]  �;  �   ��  \       ��A            � 1  �  �  +         ����  < >          � � l�       s  x<  8    ��  \       ��A            � 2  �  �  +         ����  ? A          � � s�       �  h=  �(   ��  \       ��A            � 3  �  �  +         ����  3 5          � � y�         F  ȼ   ��  ]
     	  ��B           	 � 8  �  �  ,         ����  6 7          � � ��         "G  T�   ��  ]     	  ��B           	 � 9  �  �  ,         ����  9 :          � � ��       8  0H  ��   ��  ]     	  ��B           	 � :  �  �  ,         ����  = >          � � ��       S  >I  l�   ��  ]     	  ��B           	 � ;  �  �  ,         ����  @ A          � � ��       n  LJ  ��   ��  ]     	  ��B           	 � <  �  �  ,         ����  C D          � � ��       �  ZK  ��   ��  ]     	  ��B           	 � =  �  �  ,         ����  6 7          � � ��       X	  �T  ��   ��  ^
     
  ��C           
 8  �  �  -         ����  9 :          � � ��       y	  "V  v�   ��  ^     
  ��C           
 9  �  �  -         ����  < =          � � ��       �	  NW  Z�   ��  ^     
  ��C           
 :  �  �  -         ����  @ A          � � ��       �	  zX  >�   ��  ^     
  ��C           
 ;  �  �  -         ����  C E          � ��       �	  �Y  "�   ��  ^     
  ��C           
  <  �  �  -         ����  F H          � ��       �	  �Z  �   ��  ^     
  ��C           
 � =  �  �  -         ����  9 :          � �� n     *  ^e  h�   ��  _
       ���            B  �  �  �         ����  < =          � �� o     R  �f  ��   ��  _       ���            C  �  �  �         ����  ? @          � �� p     z  �g  X�   ��  _       ���            D  �  �  �         ����  C D          � !�� q     �  <i  ��   ��  _       ���            
E  �  �  �         ����  F H          � '�� r     �  �j  H�   ��  _       ���            	F  �  �  �         ����  J K          � -�� s     �  �k  �   ��  _       ���            G  �  �  �         ����  ; =          � .�� x     �  Lw  �   ��  `
       ���            B  �  �  �         ����  > @          � 4 � y     �  �x  $!   ��  `       ���            C  �  �  �         ����  A C          � :� z     �  z  l3   ��  `       ���            D  �  �  �         ����  F H          � @� {       �{  �E   ��  `       ���            E  �  �  �         ����  J K          � F� |     >  �|  �W   ��  `       ���            F  �  �  �         ����  M O          � L � }     m  T~  Dj   ��  `       ���            G  �  �  �         ����  > ?          � L'� �     m  ��  ��   ��  a
       ��D            "L  �  �  �         ����  A C          � R/� �     �  F�  ԫ   ��  a       ��D            !M  �  �  �         ����  D F          � X7� �     �  ̍  (�   ��  a       ��D             N  �  �  �         ����  I K          � ^?� �       R�  |�   ��  a       ��D            O  �  �  �         ����  M O          dG� �     I  ؐ  ��   ��  a       ��D            P  �  �  �         ����  Q S          	jO� �     �  ^�  $   ��  a       ��D            Q  �  �  �         ����  B D          jV� �     �  ��  �[	   ��  b
       ��w            .L  �  �  
         ����  E G          p^� �     4  ^�  �t	   ��  b       ��w            -M  �  �  
         ����  I J          vf� �     s  �  �	   ��  b       ��w            ,N  �  �  
         ����  N P          #|n� �     �  ��  ��	   ��  b       ��w            +O  �  �  
         ����  R T          )�v�     �  J�  V�	   ��  b       ��w            *P  �  �  
         ����  V X          /�~�     0  �  ��	   ��  b       ��w            )Q  �  �  
         ����  E F          1���     (  :�  �c   ��  c
       ��x            ;V  �  �           ����  H J          7���     p  ��  �   ��  c       ��x            :W  �  �           ����  L M          =���     �  ��  ��   ��  c       ��x            9X  �  �           ����  Q S          C��!�        ��   �   ��  c       ��x            8Y  �  �           ����  U W          I��'�     H  B�   �   ��  c       ��x            7Z  �  �           ����  Z [          O��-�     �  �  @�   ��  c       ��x            6[  �  �           ����  2 3          x � 8j       �  h=  �(      �
     �   �            � .  �  �  �         ����  4 6          | � ?n       �  X>  1       �     �   �            � /  �  �  �         ����  7 9          � � Fr       �  H?  �9   ��  �     �   �            � 0  �  �  �         ����  ; =          � � Mv       �  8@  �A   ��  �     �   �            � 1  �  �  �         ����  > @          � � Tz       �  (A  hJ   ��  �     �   �            � 2  �  �  �         ����  A C          � � [~       �  B  �R   ��  �     �   �            � 3  �  �  �         ����  5 6          � � ay       z  �J  ��   ��  �
     �   �           	 � 8  �  �  �         ����  7 9          � � h}       �  �K  4�   ��  �     �   �           	 � 9  �  �  �         ����  : <          � � o�       �  �L  �    ��  �     �   �           	 � :  �  �  �         ����  > @          � � v�       �  �M  L   ��  �     �   �           	 � ;  �  �  �         ����  A C          � � }�       �  �N  �   ��  �     �   �           	 � <  �  �  �         ����  D F          � � ��         
P  d    ��  �     �   �           	 � =  �  �  �         ����  7 9          � � ��       �	  �Y  "�   ��  �
     �   �           
 8  �  �  �         ����  : <          � � ��       �	  �Z  �   ��  �     �   �           
 9  �  �  �         ����  = ?          � � ��       
  �[  ��   ��  �     �   �           
 :  �  �  �         ����  A C          � � ��       ?
  *]  �    ��  �     �   �           
 ;  �  �  �         ����  E F          � � ��       `
  V^  �   ��  �     �   �           
  <  �  �  �         ����  H J          � � ��       �
  �_  �   ��  �     �   �           
 � =  �  �  �         ����  : ;          � � �� n     �  j  ��   ��  �
     �   �            B  �  �  �         ����  = >          � �� o     �  Xk      ��  �     �   �            C  �  �  �         ����  @ A          � �� p     
  �l  �   ��  �     �   �            D  �  �  �         ����  D F          � �� q     2  �m  '   ��  �     �   �            
E  �  �  �         ����  H J          � �� r     Z  6o  �6   ��  �     �   �            	F  �  �  �         ����  K M          � �� s     �  �p   F   ��  �     �   �            G  �  �  �         ����  = >          � �� x       �{  �K   ��  �
     �   �            B  �  �  �         ����  @ A          � !�� y     M  d}  ^   ��  �     �   �            C  �  �  �         ����  C D          � '�� z     |  �~  \p   ��  �     �   �            D  �  �  �         ����  H I          � -�� {     �  4�  ��   ��  �     �   �            E  �  �  �         ����  K M          � 3 � |     �  ��  �   ��  �     �   �            F  �  �  �         ����  O Q          � 9� }     	  �  4�   ��  �     �   �            G  �  �  �         ����  ? A          � 9� �       p�   �   ��  �
     �   I            "L  �  �  �         ����  C D          � ?� �     L  ��  t�   ��  �     �   I            !M  �  �  �         ����  F G          � E� �     �  |�  �   ��  �     �   I             N  �  �  �         ����  K L          � K'� �     �  �     ��  �     �   I            O  �  �  �         ����  O P          � Q/� �     �  ��  p-   ��  �     �   I            P  �  �  �         ����  S T           W7� �     (  �  �B   ��  �     �   I            Q  �  �  �         ����  E F          W>� �     �  j�  6�	   ��  �
     �   �            .L  �  �           ����  H J          ]F� �     �  �  Һ	   ��  �     �   �            -M  �  �           ����  L M          cN� �     '  ��  n�	   ��  �     �   �            ,N  �  �           ����  Q S          iV� �     f  V�  
�	   ��  �     �   �            +O  �  �           ����  U W           o^� �     �  ��  �
   ��  �     �   �            *P  �  �           ����  Z [          &uf� �     �  ��  B
   ��  �     �   �            )Q  �  �           ����  H I          (~l�     �  �  ��   ��  �
     �   �            ;V  �  �           ����  K M          .�t�     0  ��  ��   ��  �     �   �            :W  �  �           ����  O P          4�|�     x  n�  ��   ��  �     �   �            9X  �  �           ����  T V          :���     �  0�      ��  �     �   �            8Y  �  �           ����  Y Z          @���       ��      ��  �     �   �            7Z  �  �           ����  ] _          F��$�     P  ��  @;   ��  �     �   �            6[  �  �           ����   9 :          � r f       �  (7  h�      m
       ��}            � .  �  �  =         ����   < =          � v j         8  ��       m       ��}            � /  �  �  =         ����   ? @          z n       #  9  H   ��  m       ��}            � 0  �  �  =         ����   C D          ~ r       9  �9  �	   ��  m       ��}            � 1  �  �  =         ����   F H          � v       O  �:  (   ��  m       ��}            � 2  �  �  =         ����   J K          #� z       e  �;  �   ��  m       ��}            � 3  �  �  =         ����   = >          $� u       �  �D  (�   ��  n
     	  ���           	 � 8  �  �  I         ����   @ A          *� y       �  �E  ��   ��  n     	  ���           	 � 9  �  �  I         ����   C D          "0� }         �F  @�   ��  n     	  ���           	 � :  �  �  I         ����   H I          (6� �       +  �G  ��   ��  n     	  ���           	 � ;  �  �  I         ����   K M          .<� �       F  �H  X�   ��  n     	  ���           	 � <  �  �  I         ����   O Q          4B� �       a  �I  ��   ��  n     	  ���           	 � =  �  �  I         ����   A B          6B� �       ,	  fS  b�   ��  o
     
  ���           
 8  �  �  U         ����   D E          <H� �       M	  �T  F�   ��  o     
  ���           
 9  �  �  U         ����   G I          BN� �       n	  �U  *�   ��  o     
  ���           
 :  �  �  U         ����   L N          HT� �       �	  �V  �   ��  o     
  ���           
 ;  �  �  U         ����   P R          NZ� �       �	  X  ��   ��  o     
  ���           
  <  �  �  U         ����   T V          T`� �       �	  BY  ��   ��  o     
  ���           
 � =  �  �  U         ����   E F          _i� � n     �  �c  ��   ��  p
       ���            B  �  �  a         ����   H J          fp� � o     "  e   �   ��  p       ���            C  �  �  a         ����   L M          mw� � p     J  bf  ��   ��  p       ���            D  �  �  a         ����   Q S          t~� � q     r  �g  �   ��  p       ���            
E  �  �  a         ����   U W          {�� � r     �  �h  ��   ��  p       ���            	F  �  �  a         ����   Z [          ��� � s     �  @j   �   ��  p       ���            G  �  �  a         ����   I J          ��� � x     N  �u  ��   ��  q
       ���            B  �  �  m         ����   M N          ��� � y     }  $w  �   ��  q       ���            C  �  �  m         ����   P R          ��� � z     �  �x     ��  q       ���            D  �  �  m         ����   V X          ��� � {     �  �y  d1   ��  q       ���            E  �  �  m         ����   Z \          ��� � |     
  \{  �C   ��  q       ���            F  �  �  m         ����   _ a          ��� � }     9  �|  �U   ��  q       ���            G  �  �  m         ����   L M          ��� � �     5  0�  ��   ��  r
       ��+            "L  �  �  �         ����   O Q          ��� � �     l  ��  ��   ��  r       ��+            !M  �  �  �         ����   S U          ��� � �     �  <�  H�   ��  r       ��+             N  �  �  �         ����   Y [          ��� � �     �    ��   ��  r       ��+            O  �  �  �         ����   ^ _          ��� � �       H�  ��   ��  r       ��+            P  �  �  �         ����   b d          ��� � �     H  ΐ  D�   ��  r       ��+            Q  �  �  �         ����   Q R          ��� � �     �  *�  vD	   ��  s
       ��=            .L  �  �  �         ����   U V          ��� � �     �  Ο  ]	   ��  s       ��=            -M  �  �  �         ����   Y [          ��� � �     7  r�  �u	   ��  s       ��=            ,N  �  �  �         ����   ` a          ��� � �     v  �  J�	   ��  s       ��=            +O  �  �  �         ����   d f          ��� �     �  ��  �	   ��  s       ��=            *P  �  �  �         ����   i k          ��� �     �  ^�  ��	   ��  s       ��=            )Q  �  �  �         ����   U V          �     �  ��  �J   ��  t
       ��>            ;V  �  �  �         ����   Y [          �     0  l�  �f   ��  t       ��>            :W  �  �  �         ����   ^ _          �     x  .�  ��   ��  t       ��>            9X  �  �  �         ����   d f           �     �  �   �   ��  t       ��>            8Y  �  �  �         ����   i k          %'&�       ��   �   ��  t       ��>            7Z  �  �  �         ����   o p          -/, �     P  t�  @�   ��  t       ��>            6[  �  �  �         ����  9 :          � � r f       �  45  ��      �
       ��            � .  �  �  ?         ����  < =          � v j       �  $6  D�       �       ��            � /  �  �  ?         ����  ? @          z n       �  7  ��   ��  �       ��            � 0  �  �  ?         ����  C D          ~ r         8  $�   ��  �       ��            � 1  �  �  ?         ����  F H          � v       "  �8  �    ��  �       ��            � 2  �  �  ?         ����  J K          � z       8  �9  	   ��  �       ��            � 3  �  �  ?         ����  = >          � u       �  �B  ��   ��  �
     	  ���           	 � 8  �  �  K         ����  @ A           � y       �  �C  ,�   ��  �     	  ���           	 � 9  �  �  K         ����  C D          "&� }       �  �D  ��   ��  �     	  ���           	 � :  �  �  K         ����  H I          (,� �       �  �E  D�   ��  �     	  ���           	 � ;  �  �  K         ����  K M          .2� �         �F  ��   ��  �     	  ���           	 � <  �  �  K         ����  O Q          48� �       /  �G  \�   ��  �     	  ���           	 � =  �  �  K         ����  A B          68� �       �  rQ  �   ��  �
     
  ���           
 8  �  �  W         ����  D E          <>� �       	  �R  ʌ   ��  �     
  ���           
 9  �  �  W         ����  G I          BD� �       7	  �S  ��   ��  �     
  ���           
 :  �  �  W         ����  L N          HJ� �       X	  �T  ��   ��  �     
  ���           
 ;  �  �  W         ����  P R          NP� �       y	  "V  v�   ��  �     
  ���           
  <  �  �  W         ����  T V          TV� �       �	  NW  Z�   ��  �     
  ���           
 � =  �  �  W         ����  E F          __� � n     �  �a  8�   ��  �
       ���            B  �  �  c         ����  H J          ff� � o     �  $c  ��   ��  �       ���            C  �  �  c         ����  L M          mm� � p       nd  (�   ��  �       ���            D  �  �  c         ����  Q S          tt� � q     6  �e  ��   ��  �       ���            
E  �  �  c         ����  U W          {{� � r     ^  g  �   ��  �       ���            	F  �  �  c         ����  Z [          ��� � s     �  Lh  ��   ��  �       ���            G  �  �  c         ����  I J          ��� � x       �s  (�   ��  �
       ���            B  �  �  o         ����  M N          ��� � y     <  0u  p�   ��  �       ���            C  �  �  o         ����  P R          ��� � z     k  �v  �   ��  �       ���            D  �  �  o         ����  V X          ��� � {     �   x      ��  �       ���            E  �  �  o         ����  Z \          ��� � |     �  hy  H*   ��  �       ���            F  �  �  o         ����  _ a          ��� � }     �  �z  �<   ��  �       ���            G  �  �  o         ����  L M          ��� � �     �  <�  He   ��  �
       ��0            "L  �  �  �         ����  O Q          ��� � �     &    �z   ��  �       ��0            !M  �  �  �         ����  S U          ��� � �     ]  H�  ��   ��  �       ��0             N  �  �  �         ����  Y [          ��� � �     �  ΋  D�   ��  �       ��0            O  �  �  �         ����  ^ _          ��� � �     �  T�  ��   ��  �       ��0            P  �  �  �         ����  b d          ��� � �       ڎ  ��   ��  �       ��0            Q  �  �  �         ����  Q R          ��� � �     n  6�  *'	   ��  �
       ��I            .L  �  �  �         ����  U V          ��� � �     �  ڝ  �?	   ��  �       ��I            -M  �  �  �         ����  Y [          ��� � �     �  ~�  bX	   ��  �       ��I            ,N  �  �  �         ����  ` a          ��� � �     +  "�  �p	   ��  �       ��I            +O  �  �  �         ����  d f          ��� �     j  Ƣ  ��	   ��  �       ��I            *P  �  �  �         ����  i k          ��� �     �  j�  6�	   ��  �       ��I            )Q  �  �  �         ����  U V          ��     �  ��  `+   ��  �
       ��J            ;V  �  �  �         ����  Y [          �     �  x�  �G   ��  �       ��J            :W  �  �  �         ����  ^ _          �     (  :�  �c   ��  �       ��J            9X  �  �  �         ����  d f           �     p  ��  �   ��  �       ��J            8Y  �  �  �         ����  i k          %&�     �  ��  ��   ��  �       ��J            7Z  �  �  �         ����  o p          -%, �        ��   �   ��  �       ��J            6[  �  �  �         ����  9 :          � r f       �  �4  P�      ;
       ��~            � .  �  �  >         ����  < =          � 
v j       �  �5  ��       ;       ��~            � /  �  �  >         ����  ? @          z n       �  �6  0�   ��  ;       ��~            � 0  �  �  >         ����  C D          ~ r         �7  ��   ��  ;       ��~            � 1  �  �  >         ����  F H          � v         �8  �   ��  ;       ��~            � 2  �  �  >         ����  J K          "� z       /  �9  �   ��  ;       ��~            � 3  �  �  >         ����  = >          #� u       �  ,B  ��   ��  <
     	  ���           	 � 8  �  �  J         ����  @ A          )� y       �  :C  D�   ��  <     	  ���           	 � 9  �  �  J         ����  C D          "/� }       �  HD  Ъ   ��  <     	  ���           	 � :  �  �  J         ����  H I          (5� �       �  VE  \�   ��  <     	  ���           	 � ;  �  �  J         ����  K M          .;� �       
  dF  �   ��  <     	  ���           	 � <  �  �  J         ����  O Q          4A� �       %  rG  t�   ��  <     	  ���           	 � =  �  �  J         ����  A B          6A� �       �  Q  �{   ��  =
     
  ���           
 8  �  �  V         ����  D E          <G� �       	  :R  ~�   ��  =     
  ���           
 9  �  �  V         ����  G I          BM� �       ,	  fS  b�   ��  =     
  ���           
 :  �  �  V         ����  L N          HS� �       M	  �T  F�   ��  =     
  ���           
 ;  �  �  V         ����  P R          NY� �       n	  �U  *�   ��  =     
  ���           
  <  �  �  V         ����  T V          T_� �       �	  �V  �   ��  =     
  ���           
 � =  �  �  V         ����  E F          _h� � n     �  va  ��   ��  >
       ���            B  �  �  b         ����  H J          fo� � o     �  �b   �   ��  >       ���            C  �  �  b         ����  L M          mv� � p       
d  x�   ��  >       ���            D  �  �  b         ����  Q S          t}� � q     *  Te  �   ��  >       ���            
E  �  �  b         ����  U W          {�� � r     R  �f  h�   ��  >       ���            	F  �  �  b         ����  Z [          ��� � s     z  �g  ��   ��  >       ���            G  �  �  b         ����  I J          ��� � x        ds  �   ��  ?
       ���            B  �  �  n         ����  M N          ��� � y     /  �t  \�   ��  ?       ���            C  �  �  n         ����  P R          ��� � z     ^  4v  �    ��  ?       ���            D  �  �  n         ����  V X          ��� � {     �  �w  �   ��  ?       ���            E  �  �  n         ����  Z \          ��� � |     �  y  4%   ��  ?       ���            F  �  �  n         ����  _ a          ��� � }     �  lz  |7   ��  ?       ���            G  �  �  n         ����  L M          ��� � �     �  ؆  �_   ��  @
       ��6            "L  �  �  �         ����  O Q          ��� � �       ^�  $u   ��  @       ��6            !M  �  �  �         ����  S U          ��� � �     O  �  x�   ��  @       ��6             N  �  �  �         ����  Y [          ��� � �     �  j�  ̟   ��  @       ��6            O  �  �  �         ����  ^ _          ��� � �     �  ��   �   ��  @       ��6            P  �  �  �         ����  b d          ��� � �     �  v�  t�   ��  @       ��6            Q  �  �  �         ����  Q R          ��� � �     _  қ  N!	   ��  A
       ��U            .L  �  �  �         ����  U V          ��� � �     �  v�  �9	   ��  A       ��U            -M  �  �  �         ����  Y [          ��� � �     �  �  �R	   ��  A       ��U            ,N  �  �  �         ����  ` a          ��� � �       ��  "k	   ��  A       ��U            +O  �  �  �         ����  d f          ��� �     [  b�  ��	   ��  A       ��U            *P  �  �  �         ����  i k          ��� �     �  �  Z�	   ��  A       ��U            )Q  �  �  �         ����  U V          �     �  R�   %   ��  B
       ��V            ;V  �  �  �         ����  Y [          �     �  �  @A   ��  B       ��V            :W  �  �  �         ����  ^ _          �       ֵ  `]   ��  B       ��V            9X  �  �  �         ����  d f           �     `  ��  �y   ��  B       ��V            8Y  �  �  �         ����  i k          %&&�     �  Z�  ��   ��  B       ��V            7Z  �  �  �         ����  o p          -., �     �  �  ��   ��  B       ��V            6[  �  �  �         ����  9 :          � � r f       c  �;  �      �
       ���            � .  �  �  @         ����  < =          � � v j       y  �<  #       �       ���            � /  �  �  @         ����  ? @          z n       �  �=  x+   ��  �       ���            � 0  �  �  @         ����  C D          
~ r       �  �>  �3   ��  �       ���            � 1  �  �  @         ����  F H          � v       �  �?  X<   ��  �       ���            � 2  �  �  @         ����  J K          � z       �  �@  �D   ��  �       ���            � 3  �  �  @         ����  ; =          � u       R  4I  �   ��  �
     	  ���           	 � 8  �  �  L         ����  > @          � y       m  BJ  ��   ��  �     	  ���           	 � 9  �  �  L         ����  A C          "#� }       �  PK   �   ��  �     	  ���           	 � :  �  �  L         ����  F H          ()� �       �  ^L  ��   ��  �     	  ���           	 � ;  �  �  L         ����  J K          ./� �       �  lM  8   ��  �     	  ���           	 � <  �  �  L         ����  M O          45� �       �  zN  �   ��  �     	  ���           	 � =  �  �  L         ����  A B          65� �       �	  X  ��   ��  �
     
  ���           
 8  �  �  X         ����  D E          <;� �       �	  BY  ��   ��  �     
  ���           
 9  �  �  X         ����  G I          BA� �       �	  nZ  ��   ��  �     
  ���           
 :  �  �  X         ����  L N          HG� �       
  �[  ��   ��  �     
  ���           
 ;  �  �  X         ����  P R          NM� �       4
  �\  ��   ��  �     
  ���           
  <  �  �  X         ����  T V          TS� �       U
  �]  f	   ��  �     
  ���           
 � =  �  �  X         ����  E F          _\� � n     �  ~h  ��   ��  �
       ���            B  �  �  d         ����  H J          fc� � o     �  �i  `�   ��  �       ���            C  �  �  d         ����  L M          mj� � p     �  k  �   ��  �       ���            D  �  �  d         ����  Q S          tq� � q       \l  P   ��  �       ���            
E  �  �  d         ����  U W          {x� � r     *  �m  �#   ��  �       ���            	F  �  �  d         ����  Z [          �� � s     R  �n  @3   ��  �       ���            G  �  �  d         ����  I J          ��� � x     �  lz  |7   ��  �
       ���            B  �  �  p         ����  M N          ��� � y       �{  �I   ��  �       ���            C  �  �  p         ����  P R          ��� � z     H  <}  \   ��  �       ���            D  �  �  p         ����  V X          ��� � {     w  �~  Tn   ��  �       ���            E  �  �  p         ����  Z \          ��� � |     �  �  ��   ��  �       ���            F  �  �  p         ����  _ a          ��� � }     �  t�  �   ��  �       ���            G  �  �  p         ����  L M          ��� � �     �  ��  @�   ��  �
       ��;            "L  �  �  �         ����  O Q          ��� � �       f�  ��   ��  �       ��;            !M  �  �  �         ����  S U          ��� � �     K  �  ��   ��  �       ��;             N  �  �  �         ����  Y [          ��� � �     �  r�  <   ��  �       ��;            O  �  �  �         ����  ^ _          ��� � �     �  ��  �   ��  �       ��;            P  �  �  �         ����  b d          ��� � �     �  ~�  �,   ��  �       ��;            Q  �  �  �         ����  Q R          ��� � �     m  ڢ  Ɗ	   ��  �
       ��a            .L  �  �  �         ����  U V          ��� � �     �  ~�  b�	   ��  �       ��a            -M  �  �  �         ����  Y [          ��� � �     �  "�  ��	   ��  �       ��a            ,N  �  �  �         ����  ` a          ��� � �     *  Ƨ  ��	   ��  �       ��a            +O  �  �  �         ����  d f          ��� �     i  j�  6�	   ��  �       ��a            *P  �  �  �         ����  i k          ��� �     �  �  �
   ��  �       ��a            )Q  �  �  �         ����  U V          ��     �  Z�  ��   ��  �
       ��b            ;V  �  �  �         ����  Y [          �     �  �  ��   ��  �       ��b            :W  �  �  �         ����  ^ _          
�     8  ޼  ��   ��  �       ��b            9X  �  �  �         ����  d f           �     �  ��   �   ��  �       ��b            8Y  �  �  �         ����  i k          %&�     �  b�      ��  �       ��b            7Z  �  �  �         ����  o p          -", �       $�  @"   ��  �       ��b            6[  �  �  �         ����  ; =          � r f       ?  H:  �      
       ���            � .  �  �  B         ����  > @          � v j       U  8;  �              ���            � /  �  �  B         ����  A C          z n       k  (<  h   ��         ���            � 0  �  �  B         ����  F H          !~ r       �  =  �%   ��         ���            � 1  �  �  B         ����  J K          '� v       �  >  H.   ��         ���            � 2  �  �  B         ����  M O          -� z       �  �>  �6   ��         ���            � 3  �  �  B         ����  ? A          .� u       *  �G  h�   ��  
       ���           	 � 8  �  �  N         ����  C D          4� y       E  �H  ��   ��         ���           	 � 9  �  �  N         ����  F G          ":� }       `  �I  ��   ��         ���           	 � :  �  �  N         ����  K L          (@� �       {  �J  �   ��         ���           	 � ;  �  �  N         ����  O P          .F� �       �  �K  ��   ��         ���           	 � <  �  �  N         ����  S T          4L� �       �  �L  $   ��         ���           	 � =  �  �  N         ����  B D          6L� �       �	  �V  ·   ��  	
     	  ���           
 8  �  �  Z         ����  E G          <R� �       �	  �W  ��   ��  	     	  ���           
 9  �  �  Z         ����  I J          BX� �       �	  �X  ��   ��  	     	  ���           
 :  �  �  Z         ����  N P          H^� �       �	  
Z  n�   ��  	     	  ���           
 ;  �  �  Z         ����  R T          Nd� �       
  6[  R�   ��  	     	  ���           
  <  �  �  Z         ����  V X          Tj� �       )
  b\  6�   ��  	     	  ���           
 � =  �  �  Z         ����  F H          _s� � n     Z  �f  (�   ��  

     
  ���            B  �  �  f         ����  J K          fz� � o     �  8h  ��   ��  
     
  ���            C  �  �  f         ����  M O          m�� � p     �  �i  �   ��  
     
  ���            D  �  �  f         ����  S T          t�� � q     �  �j  �   ��  
     
  ���            
E  �  �  f         ����  W Y          {�� � r     �  l     ��  
     
  ���            	F  �  �  f         ����  [ ]          ��� � s     "  `m  �    ��  
     
  ���            G  �  �  f         ����  J L          ��� � x     �  �x  ,#   ��  
       ���            B  �  �  r         ����  N O          ��� � y     �  Dz  t5   ��         ���            C  �  �  r         ����  R S          ��� � z       �{  �G   ��         ���            D  �  �  r         ����  X Y          ��� � {     C  }  Z   ��         ���            E  �  �  r         ����  \ ^          ��� � |     r  |~  Ll   ��         ���            F  �  �  r         ����  a b          ��� � }     �  �  �~   ��         ���            G  �  �  r         ����  N P          ��� � �     �  P�  `�   ��  
       ��@            "L  �  �  �         ����  R T          ��� � �     �  ֍  ��   ��         ��@            !M  �  �  �         ����  V X          ��� � �       \�  �   ��         ��@             N  �  �  �         ����  \ ^          ��� � �     J  �  \�   ��         ��@            O  �  �  �         ����  a c          ��� � �     �  h�  �   ��         ��@            P  �  �  �         ����  f h          ��� � �     �  �     ��         ��@            Q  �  �  �         ����  T U          ��� � �     1  J�  Vs	   ��  
       ��m            .L  �  �            ����  X Y          ��� � �     p  �  �	   ��         ��m            -M  �  �            ����  \ ^          ��� � �     �  ��  ��	   ��         ��m            ,N  �  �            ����  c d          ��� � �     �  6�  *�	   ��         ��m            +O  �  �            ����  h i          ��� �     -  ڧ  ��	   ��         ��m            *P  �  �            ����  m o          �� �     l  ~�  b�	   ��         ��m            )Q  �  �            ����  V X          �     h  ʷ  �|   ��  
       ��n            ;V  �  �           ����  [ \          �     �  ��  ��   ��         ��n            :W  �  �           ����  _ a          !�     �  N�  �   ��         ��n            9X  �  �           ����  f h          ) �     @  �   �   ��         ��n            8Y  �  �           ����  k m          %1&�     �  Ҿ   �   ��         ��n            7Z  �  �           ����  p r          -9, �     �  ��  @	   ��         ��n            6[  �  �           ����  : ;          � � r f         �8  x�      m
       ���            � .  �  �  A         ����  = >          � v j       1  �9  �       m       ���            � /  �  �  A         ����  @ A          z n       G  �:  X   ��  m       ���            � 0  �  �  A         ����  D F          ~ r       ]  �;  �   ��  m       ���            � 1  �  �  A         ����  H J          � v       s  x<  8    ��  m       ���            � 2  �  �  A         ����  K M          � z       �  h=  �(   ��  m       ���            � 3  �  �  A         ����  > ?          � u         F  ȼ   ��  n
     	  ���           	 � 8  �  �  M         ����  A C          !� y         "G  T�   ��  n     	  ���           	 � 9  �  �  M         ����  D F          "'� }       8  0H  ��   ��  n     	  ���           	 � :  �  �  M         ����  I K          (-� �       S  >I  l�   ��  n     	  ���           	 � ;  �  �  M         ����  M O          .3� �       n  LJ  ��   ��  n     	  ���           	 � <  �  �  M         ����  Q S          49� �       �  ZK  ��   ��  n     	  ���           	 � =  �  �  M         ����  B D          69� �       X	  �T  ��   ��  o
     
  ���           
 8  �  �  Y         ����  E G          <?� �       y	  "V  v�   ��  o     
  ���           
 9  �  �  Y         ����  I J          BE� �       �	  NW  Z�   ��  o     
  ���           
 :  �  �  Y         ����  N P          HK� �       �	  zX  >�   ��  o     
  ���           
 ;  �  �  Y         ����  R T          NQ� �       �	  �Y  "�   ��  o     
  ���           
  <  �  �  Y         ����  V X          TW� �       �	  �Z  �   ��  o     
  ���           
 � =  �  �  Y         ����  F H          _`� � n     *  ^e  h�   ��  p
       ���            B  �  �  e         ����  J K          fg� � o     R  �f  ��   ��  p       ���            C  �  �  e         ����  M O          mn� � p     z  �g  X�   ��  p       ���            D  �  �  e         ����  S T          tu� � q     �  <i  ��   ��  p       ���            
E  �  �  e         ����  W Y          {|� � r     �  �j  H�   ��  p       ���            	F  �  �  e         ����  [ ]          ��� � s     �  �k  �   ��  p       ���            G  �  �  e         ����  I J          ��� � x     �  Lw  �   ��  q
       ���            B  �  �  q         ����  M N          ��� � y     �  �x  $!   ��  q       ���            C  �  �  q         ����  P R          ��� � z     �  z  l3   ��  q       ���            D  �  �  q         ����  V X          ��� � {       �{  �E   ��  q       ���            E  �  �  q         ����  Z \          ��� � |     >  �|  �W   ��  q       ���            F  �  �  q         ����  _ a          ��� � }     m  T~  Dj   ��  q       ���            G  �  �  q         ����  M N          ��� � �     m  ��  ��   ��  r
       ��E            "L  �  �  �         ����  Q R          ��� � �     �  F�  ԫ   ��  r       ��E            !M  �  �  �         ����  U V          ��� � �     �  ̍  (�   ��  r       ��E             N  �  �  �         ����  [ \          ��� � �       R�  |�   ��  r       ��E            O  �  �  �         ����  _ a          ��� � �     I  ؐ  ��   ��  r       ��E            P  �  �  �         ����  d f          ��� � �     �  ^�  $   ��  r       ��E            Q  �  �  �         ����  R T          ��� � �     �  ��  �[	   ��  s
       ��y            .L  �  �           ����  V X          ��� � �     4  ^�  �t	   ��  s       ��y            -M  �  �           ����  [ \          ��� � �     s  �  �	   ��  s       ��y            ,N  �  �           ����  a c          ��� � �     �  ��  ��	   ��  s       ��y            +O  �  �           ����  f h          ��� �     �  J�  V�	   ��  s       ��y            *P  �  �           ����  k m          ��� �     0  �  ��	   ��  s       ��y            )Q  �  �           ����  V X          ��     (  :�  �c   ��  t
       ��z            ;V  �  �           ����  [ \          �     p  ��  �   ��  t       ��z            :W  �  �           ����  _ a          �     �  ��  ��   ��  t       ��z            9X  �  �           ����  f h           �        ��   �   ��  t       ��z            8Y  �  �           ����  k m          %&�     H  B�   �   ��  t       ��z            7Z  �  �           ����  p r          -&, �     �  �  @�   ��  t       ��z            6[  �  �           ����    9 :          | � Bf       �  (7  h�      
       ��^            � .  �  �  
         ����    < =          � � Ij         8  ��              ��^            � /  �  �  
         ����    ? @          � � Pn       #  9  H   ��         ��^            � 0  �  �  
         ����    C D          � � Wr       9  �9  �	   ��         ��^            � 1  �  �  
         ����    F H          � � ^v       O  �:  (   ��         ��^            � 2  �  �  
         ����    J K          � � ez       e  �;  �   ��         ��^            � 3  �  �  
         ����    = >          � � ku       �  �D  (�   ��  �
     	  ��_           	 � 8  �  �           ����    @ A          � � ry       �  �E  ��   ��  �     	  ��_           	 � 9  �  �           ����    C D          � � y}         �F  @�   ��  �     	  ��_           	 � :  �  �           ����    H I          � � ��       +  �G  ��   ��  �     	  ��_           	 � ;  �  �           ����    K M          � � ��       F  �H  X�   ��  �     	  ��_           	 � <  �  �           ����    O Q          � � ��       a  �I  ��   ��  �     	  ��_           	 � =  �  �           ����    ? A          � � ��       ,	  fS  b�   ��  �
     
  ��`           
 8  �  �           ����    C D          � � ��       M	  �T  F�   ��  �     
  ��`           
 9  �  �           ����    F G          � � ��       n	  �U  *�   ��  �     
  ��`           
 :  �  �           ����    K L          � � ��       �	  �V  �   ��  �     
  ��`           
 ;  �  �           ����    O P          � � ��       �	  X  ��   ��  �     
  ��`           
  <  �  �           ����    S T          � � ��       �	  BY  ��   ��  �     
  ��`           
 � =  �  �           ����    D E          � �� n     �  �c  ��   ��  �
       ��a            B  �  �           ����    G H          � �� o     "  e   �   ��  �       ��a            C  �  �           ����    J L          � �� p     J  bf  ��   ��  �       ��a            D  �  �           ����    P Q          � �� q     r  �g  �   ��  �       ��a            
E  �  �           ����    T U          � �� r     �  �h  ��   ��  �       ��a            	F  �  �           ����    X Z          �  �� s     �  @j   �   ��  �       ��a            G  �  �           ����    H I          � !�� x     N  �u  ��   ��  �
       ��b            B  �  �           ����    K M          � '�� y     }  $w  �   ��  �       ��b            C  �  �           ����    O P          � -�� z     �  �x     ��  �       ��b            D  �  �           ����    T V          � 3� {     �  �y  d1   ��  �       ��b            E  �  �           ����    Y Z          � 9
� |     
  \{  �C   ��  �       ��b            F  �  �           ����    ] _          � ?� }     9  �|  �U   ��  �       ��b            G  �  �           ����    L M          � ?� �     5  0�  ��   ��  �
       ��c            "L  �  �           ����    O Q          � E!� �     l  ��  ��   ��  �       ��c            !M  �  �           ����    S U          � K)� �     �  <�  H�   ��  �       ��c             N  �  �           ����    Y [          � Q1� �     �    ��   ��  �       ��c            O  �  �           ����    ^ _          � W9� �       H�  ��   ��  �       ��c            P  �  �           ����    b d          ]A� �     H  ΐ  D�   ��  �       ��c            Q  �  �           ����    Q R          ]H� �     �  *�  vD	   ��  �
       ��?            .L  �  �  �         ����    U V          cP� �     �  Ο  ]	   ��  �       ��?            -M  �  �  �         ����    Y [          iX� �     7  r�  �u	   ��  �       ��?            ,N  �  �  �         ����    ` a          o`� �     v  �  J�	   ��  �       ��?            +O  �  �  �         ����    d f          $uh� �     �  ��  �	   ��  �       ��?            *P  �  �  �         ����    i k          *{p� �     �  ^�  ��	   ��  �       ��?            )Q  �  �  �         ����    T U          ,�v�     �  ��  �J   ��  �
       ��@            ;V  �  �  �         ����    X Y          2�~�     0  l�  �f   ��  �       ��@            :W  �  �  �         ����    \ ^          8���     x  .�  ��   ��  �       ��@            9X  �  �  �         ����    c d          >���     �  �   �   ��  �       ��@            8Y  �  �  �         ����    h i          D���       ��   �   ��  �       ��@            7Z  �  �  �         ����    m o          J�� �     P  t�  @�   ��  �       ��@            6[  �  �  �         ����   7 9          | � 6f       �  45  ��      �
       ��k            � .  �  �           ����   : <          � � =j       �  $6  D�       �       ��k            � /  �  �           ����   = ?          � � Dn       �  7  ��   ��  �       ��k            � 0  �  �           ����   A C          � � Kr         8  $�   ��  �       ��k            � 1  �  �           ����   E F          � � Rv       "  �8  �    ��  �       ��k            � 2  �  �           ����   H J          � � Yz       8  �9  	   ��  �       ��k            � 3  �  �           ����   ; =          � � _u       �  �B  ��   ��  �
     	  ��l           	 � 8  �  �           ����   > @          � � fy       �  �C  ,�   ��  �     	  ��l           	 � 9  �  �           ����   A C          � � m}       �  �D  ��   ��  �     	  ��l           	 � :  �  �           ����   F H          � � t�       �  �E  D�   ��  �     	  ��l           	 � ;  �  �           ����   J K          � � {�         �F  ��   ��  �     	  ��l           	 � <  �  �           ����   M O          � � ��       /  �G  \�   ��  �     	  ��l           	 � =  �  �           ����   ? A          � � ��       �  rQ  �   ��  �
     
  ��m           
 8  �  �           ����   C D          � � ��       	  �R  ʌ   ��  �     
  ��m           
 9  �  �           ����   F G          � � ��       7	  �S  ��   ��  �     
  ��m           
 :  �  �           ����   K L          � � ��       X	  �T  ��   ��  �     
  ��m           
 ;  �  �           ����   O P          � � ��       y	  "V  v�   ��  �     
  ��m           
  <  �  �           ����   S T          � � ��       �	  NW  Z�   ��  �     
  ��m           
 � =  �  �           ����   B D          � �� n     �  �a  8�   ��  �
       ��n            B  �  �           ����   E G          � �� o     �  $c  ��   ��  �       ��n            C  �  �           ����   I J          � �� p       nd  (�   ��  �       ��n            D  �  �           ����   N P          � �� q     6  �e  ��   ��  �       ��n            
E  �  �           ����   R T          � �� r     ^  g  �   ��  �       ��n            	F  �  �           ����   V X          �  �� s     �  Lh  ��   ��  �       ��n            G  �  �           ����   F H          � !�� x       �s  (�   ��  �
       ��o            B  �  �           ����   J K          � '�� y     <  0u  p�   ��  �       ��o            C  �  �           ����   M O          � -�� z     k  �v  �   ��  �       ��o            D  �  �           ����   S T          � 3�� {     �   x      ��  �       ��o            E  �  �           ����   W Y          � 9�� |     �  hy  H*   ��  �       ��o            F  �  �           ����   [ ]          � ?� }     �  �z  �<   ��  �       ��o            G  �  �           ����   J L          � ?� �     �  <�  He   ��  �
       ��p            "L  �  �           ����   N O          � E� �     &    �z   ��  �       ��p            !M  �  �           ����   R S          � K� �     ]  H�  ��   ��  �       ��p             N  �  �           ����   X Y          � Q%� �     �  ΋  D�   ��  �       ��p            O  �  �           ����   \ ^          � W-� �     �  T�  ��   ��  �       ��p            P  �  �           ����   a b          ]5� �       ڎ  ��   ��  �       ��p            Q  �  �           ����   P Q          ]<� �     n  6�  *'	   ��  �
       ��K            .L  �  �  �         ����   T U          cD� �     �  ڝ  �?	   ��  �       ��K            -M  �  �  �         ����   X Y          iL� �     �  ~�  bX	   ��  �       ��K            ,N  �  �  �         ����   ^ `          oT� �     +  "�  �p	   ��  �       ��K            +O  �  �  �         ����   c d          $u\� �     j  Ƣ  ��	   ��  �       ��K            *P  �  �  �         ����   h i          *{d� �     �  j�  6�	   ��  �       ��K            )Q  �  �  �         ����   T U          ,�j�     �  ��  `+   ��  �
       ��L            ;V  �  �  �         ����   X Y          2�r�     �  x�  �G   ��  �       ��L            :W  �  �  �         ����   \ ^          8�z�     (  :�  �c   ��  �       ��L            9X  �  �  �         ����   c d          >���     p  ��  �   ��  �       ��L            8Y  �  �  �         ����   h i          D���     �  ��  ��   ��  �       ��L            7Z  �  �  �         ����   m o          J�� �        ��   �   ��  �       ��L            6[  �  �  �         ����   7 9          | � >f       �  �4  P�      L
       ��x            � .  �  �  $         ����   : <          � � Ej       �  �5  ��       L       ��x            � /  �  �  $         ����   = ?          � � Ln       �  �6  0�   ��  L       ��x            � 0  �  �  $         ����   A C          � � Sr         �7  ��   ��  L       ��x            � 1  �  �  $         ����   E F          � � Zv         �8  �   ��  L       ��x            � 2  �  �  $         ����   H J          � � az       /  �9  �   ��  L       ��x            � 3  �  �  $         ����   ; =          � � gu       �  ,B  ��   ��  M
     	  ��y           	 � 8  �  �  %         ����   > @          � � ny       �  :C  D�   ��  M     	  ��y           	 � 9  �  �  %         ����   A C          � � u}       �  HD  Ъ   ��  M     	  ��y           	 � :  �  �  %         ����   F H          � � |�       �  VE  \�   ��  M     	  ��y           	 � ;  �  �  %         ����   J K          � � ��       
  dF  �   ��  M     	  ��y           	 � <  �  �  %         ����   M O          � � ��       %  rG  t�   ��  M     	  ��y           	 � =  �  �  %         ����   ? A          � � ��       �  Q  �{   ��  N
     
  ��z           
 8  �  �  &         ����   C D          � � ��       	  :R  ~�   ��  N     
  ��z           
 9  �  �  &         ����   F G          � � ��       ,	  fS  b�   ��  N     
  ��z           
 :  �  �  &         ����   K L          � � ��       M	  �T  F�   ��  N     
  ��z           
 ;  �  �  &         ����   O P          � � ��       n	  �U  *�   ��  N     
  ��z           
  <  �  �  &         ����   S T          � � ��       �	  �V  �   ��  N     
  ��z           
 � =  �  �  &         ����   B D          � �� n     �  va  ��   ��  O
       ��{            B  �  �  '         ����   E G          � �� o     �  �b   �   ��  O       ��{            C  �  �  '         ����   I J          � �� p       
d  x�   ��  O       ��{            D  �  �  '         ����   N P          � �� q     *  Te  �   ��  O       ��{            
E  �  �  '         ����   R T          � �� r     R  �f  h�   ��  O       ��{            	F  �  �  '         ����   V X          �  �� s     z  �g  ��   ��  O       ��{            G  �  �  '         ����   F H          � !�� x        ds  �   ��  P
       ��|            B  �  �  (         ����   J K          � '�� y     /  �t  \�   ��  P       ��|            C  �  �  (         ����   M O          � -�� z     ^  4v  �    ��  P       ��|            D  �  �  (         ����   S T          � 3�� {     �  �w  �   ��  P       ��|            E  �  �  (         ����   W Y          � 9� |     �  y  4%   ��  P       ��|            F  �  �  (         ����   [ ]          � ?� }     �  lz  |7   ��  P       ��|            G  �  �  (         ����   J L          � ?� �     �  ؆  �_   ��  Q
       ��}            "L  �  �  )         ����   N O          � E� �       ^�  $u   ��  Q       ��}            !M  �  �  )         ����   R S          � K%� �     O  �  x�   ��  Q       ��}             N  �  �  )         ����   X Y          � Q-� �     �  j�  ̟   ��  Q       ��}            O  �  �  )         ����   \ ^          � W5� �     �  ��   �   ��  Q       ��}            P  �  �  )         ����   a b          ]=� �     �  v�  t�   ��  Q       ��}            Q  �  �  )         ����   P Q          ]D� �     _  қ  N!	   ��  R
       ��W            .L  �  �  �         ����   T U          cL� �     �  v�  �9	   ��  R       ��W            -M  �  �  �         ����   X Y          iT� �     �  �  �R	   ��  R       ��W            ,N  �  �  �         ����   ^ `          o\� �       ��  "k	   ��  R       ��W            +O  �  �  �         ����   c d          $ud� �     [  b�  ��	   ��  R       ��W            *P  �  �  �         ����   h i          *{l� �     �  �  Z�	   ��  R       ��W            )Q  �  �  �         ����   T U          ,�r�     �  R�   %   ��  S
       ��X            ;V  �  �  �         ����   X Y          2�z�     �  �  @A   ��  S       ��X            :W  �  �  �         ����   \ ^          8���       ֵ  `]   ��  S       ��X            9X  �  �  �         ����   c d          >���     `  ��  �y   ��  S       ��X            8Y  �  �  �         ����   h i          D���     �  Z�  ��   ��  S       ��X            7Z  �  �  �         ����   m o          J�� �     �  �  ��   ��  S       ��X            6[  �  �  �         ����   7 9          | � 2f       c  �;  �      �
       ���            � .  �  �  1         ����   : <          � � 9j       y  �<  #       �       ���            � /  �  �  1         ����   = ?          � � @n       �  �=  x+   ��  �       ���            � 0  �  �  1         ����   A C          � � Gr       �  �>  �3   ��  �       ���            � 1  �  �  1         ����   E F          � � Nv       �  �?  X<   ��  �       ���            � 2  �  �  1         ����   H J          � � Uz       �  �@  �D   ��  �       ���            � 3  �  �  1         ����   ; =          � � [u       R  4I  �   ��  �
     	  ���           	 � 8  �  �  2         ����   > @          � � by       m  BJ  ��   ��  �     	  ���           	 � 9  �  �  2         ����   A C          � � i}       �  PK   �   ��  �     	  ���           	 � :  �  �  2         ����   F H          � � p�       �  ^L  ��   ��  �     	  ���           	 � ;  �  �  2         ����   J K          � � w�       �  lM  8   ��  �     	  ���           	 � <  �  �  2         ����   M O          � � ~�       �  zN  �   ��  �     	  ���           	 � =  �  �  2         ����   ? A          � � ��       �	  X  ��   ��  �
     
  ���           
 8  �  �  3         ����   C D          � � ��       �	  BY  ��   ��  �     
  ���           
 9  �  �  3         ����   F G          � � ��       �	  nZ  ��   ��  �     
  ���           
 :  �  �  3         ����   K L          � � ��       
  �[  ��   ��  �     
  ���           
 ;  �  �  3         ����   O P          � � ��       4
  �\  ��   ��  �     
  ���           
  <  �  �  3         ����   S T          � � ��       U
  �]  f	   ��  �     
  ���           
 � =  �  �  3         ����   B D          � �� n     �  ~h  ��   ��  �
       ���            B  �  �  4         ����   E G          � �� o     �  �i  `�   ��  �       ���            C  �  �  4         ����   I J          � �� p     �  k  �   ��  �       ���            D  �  �  4         ����   N P          � �� q       \l  P   ��  �       ���            
E  �  �  4         ����   R T          � �� r     *  �m  �#   ��  �       ���            	F  �  �  4         ����   V X          �  �� s     R  �n  @3   ��  �       ���            G  �  �  4         ����   F H          � !�� x     �  lz  |7   ��  �
       ���            B  �  �  5         ����   J K          � '�� y       �{  �I   ��  �       ���            C  �  �  5         ����   M O          � -�� z     H  <}  \   ��  �       ���            D  �  �  5         ����   S T          � 3�� {     w  �~  Tn   ��  �       ���            E  �  �  5         ����   W Y          � 9�� |     �  �  ��   ��  �       ���            F  �  �  5         ����   [ ]          � ?� }     �  t�  �   ��  �       ���            G  �  �  5         ����   J L          � ?	� �     �  ��  @�   ��  �
       ���            "L  �  �  6         ����   N O          � E� �       f�  ��   ��  �       ���            !M  �  �  6         ����   R S          � K� �     K  �  ��   ��  �       ���             N  �  �  6         ����   X Y          � Q!� �     �  r�  <   ��  �       ���            O  �  �  6         ����   \ ^          � W)� �     �  ��  �   ��  �       ���            P  �  �  6         ����   a b          ]1� �     �  ~�  �,   ��  �       ���            Q  �  �  6         ����   P Q          ]8� �     m  ڢ  Ɗ	   ��  �
       ��c            .L  �  �  �         ����   T U          c@� �     �  ~�  b�	   ��  �       ��c            -M  �  �  �         ����   X Y          iH� �     �  "�  ��	   ��  �       ��c            ,N  �  �  �         ����   ^ `          oP� �     *  Ƨ  ��	   ��  �       ��c            +O  �  �  �         ����   c d          $uX� �     i  j�  6�	   ��  �       ��c            *P  �  �  �         ����   h i          *{`� �     �  �  �
   ��  �       ��c            )Q  �  �  �         ����   T U          ,�f�     �  Z�  ��   ��  �
       ��d            ;V  �  �  �         ����   X Y          2�n�     �  �  ��   ��  �       ��d            :W  �  �  �         ����   \ ^          8�v�     8  ޼  ��   ��  �       ��d            9X  �  �  �         ����   c d          >�~�     �  ��   �   ��  �       ��d            8Y  �  �  �         ����   h i          D���     �  b�      ��  �       ��d            7Z  �  �  �         ����   m o          J�� �       $�  @"   ��  �       ��d            6[  �  �  �         ����   9 :          | � Jf       ?  H:  �      
       ���            � .  �  �  >         ����   < =          � � Qj       U  8;  �              ���            � /  �  �  >         ����   ? @          � � Xn       k  (<  h   ��         ���            � 0  �  �  >         ����   C D          � � _r       �  =  �%   ��         ���            � 1  �  �  >         ����   F H          � � fv       �  >  H.   ��         ���            � 2  �  �  >         ����   J K          � � mz       �  �>  �6   ��         ���            � 3  �  �  >         ����   = >          � � su       *  �G  h�   ��  
       ���           	 � 8  �  �  ?         ����   @ A          � � zy       E  �H  ��   ��         ���           	 � 9  �  �  ?         ����   C D          � � �}       `  �I  ��   ��         ���           	 � :  �  �  ?         ����   H I          � � ��       {  �J  �   ��         ���           	 � ;  �  �  ?         ����   K M          � � ��       �  �K  ��   ��         ���           	 � <  �  �  ?         ����   O Q          � � ��       �  �L  $   ��         ���           	 � =  �  �  ?         ����   ? A          � � ��       �	  �V  ·   ��  
     	  ���           
 8  �  �  @         ����   C D          � � ��       �	  �W  ��   ��       	  ���           
 9  �  �  @         ����   F G          � � ��       �	  �X  ��   ��       	  ���           
 :  �  �  @         ����   K L          � � ��       �	  
Z  n�   ��       	  ���           
 ;  �  �  @         ����   O P          � � ��       
  6[  R�   ��       	  ���           
  <  �  �  @         ����   S T          � � ��       )
  b\  6�   ��       	  ���           
 � =  �  �  @         ����   D E          � �� n     Z  �f  (�   ��  
     
  ���            B  �  �  A         ����   G H          � �� o     �  8h  ��   ��       
  ���            C  �  �  A         ����   J L          � �� p     �  �i  �   ��       
  ���            D  �  �  A         ����   P Q          � �� q     �  �j  �   ��       
  ���            
E  �  �  A         ����   T U          � �� r     �  l     ��       
  ���            	F  �  �  A         ����   X Z          �  �� s     "  `m  �    ��       
  ���            G  �  �  A         ����   H I          � !�� x     �  �x  ,#   ��  
       ���            B  �  �  B         ����   K M          � '�� y     �  Dz  t5   ��         ���            C  �  �  B         ����   O P          � -� z       �{  �G   ��         ���            D  �  �  B         ����   T V          � 3
� {     C  }  Z   ��         ���            E  �  �  B         ����   Y Z          � 9� |     r  |~  Ll   ��         ���            F  �  �  B         ����   ] _          � ?� }     �  �  �~   ��         ���            G  �  �  B         ����   L M          � ?!� �     �  P�  `�   ��  
       ���            "L  �  �  C         ����   O Q          � E)� �     �  ֍  ��   ��         ���            !M  �  �  C         ����   S U          � K1� �       \�  �   ��         ���             N  �  �  C         ����   Y [          � Q9� �     J  �  \�   ��         ���            O  �  �  C         ����   ^ _          � WA� �     �  h�  �   ��         ���            P  �  �  C         ����   b d          ]I� �     �  �     ��         ���            Q  �  �  C         ����   Q R          ]P� �     1  J�  Vs	   ��  
       ��o            .L  �  �           ����   U V          cX� �     p  �  �	   ��         ��o            -M  �  �           ����   Y [          i`� �     �  ��  ��	   ��         ��o            ,N  �  �           ����   ` a          oh� �     �  6�  *�	   ��         ��o            +O  �  �           ����   d f          $up� �     -  ڧ  ��	   ��         ��o            *P  �  �           ����   i k          *{x� �     l  ~�  b�	   ��         ��o            )Q  �  �           ����   T U          ,�~�     h  ʷ  �|   ��  
       ��p            ;V  �  �           ����   X Y          2���     �  ��  ��   ��         ��p            :W  �  �           ����   \ ^          8���     �  N�  �   ��         ��p            9X  �  �           ����   c d          >���     @  �   �   ��         ��p            8Y  �  �           ����   h i          D���     �  Ҿ   �   ��         ��p            7Z  �  �           ����   m o          J�� �     �  ��  @	   ��         ��p            6[  �  �           ����   7 9          | � :f         �8  x�      ~
       ���            � .  �  �  K         ����   : <          � � Aj       1  �9  �       ~       ���            � /  �  �  K         ����   = ?          � � Hn       G  �:  X   ��  ~       ���            � 0  �  �  K         ����   A C          � � Or       ]  �;  �   ��  ~       ���            � 1  �  �  K         ����   E F          � � Vv       s  x<  8    ��  ~       ���            � 2  �  �  K         ����   H J          � � ]z       �  h=  �(   ��  ~       ���            � 3  �  �  K         ����   ; =          � � cu         F  ȼ   ��  
     	  ���           	 � 8  �  �  L         ����   > @          � � jy         "G  T�   ��       	  ���           	 � 9  �  �  L         ����   A C          � � q}       8  0H  ��   ��       	  ���           	 � :  �  �  L         ����   F H          � � x�       S  >I  l�   ��       	  ���           	 � ;  �  �  L         ����   J K          � � �       n  LJ  ��   ��       	  ���           	 � <  �  �  L         ����   M O          � � ��       �  ZK  ��   ��       	  ���           	 � =  �  �  L         ����   ? A          � � ��       X	  �T  ��   ��  �
     
  ���           
 8  �  �  M         ����   C D          � � ��       y	  "V  v�   ��  �     
  ���           
 9  �  �  M         ����   F G          � � ��       �	  NW  Z�   ��  �     
  ���           
 :  �  �  M         ����   K L          � � ��       �	  zX  >�   ��  �     
  ���           
 ;  �  �  M         ����   O P          � � ��       �	  �Y  "�   ��  �     
  ���           
  <  �  �  M         ����   S T          � � ��       �	  �Z  �   ��  �     
  ���           
 � =  �  �  M         ����   B D          � �� n     *  ^e  h�   ��  �
       ���            B  �  �  N         ����   E G          � �� o     R  �f  ��   ��  �       ���            C  �  �  N         ����   I J          � �� p     z  �g  X�   ��  �       ���            D  �  �  N         ����   N P          � �� q     �  <i  ��   ��  �       ���            
E  �  �  N         ����   R T          � �� r     �  �j  H�   ��  �       ���            	F  �  �  N         ����   V X          �  �� s     �  �k  �   ��  �       ���            G  �  �  N         ����   F H          � !�� x     �  Lw  �   ��  �
       ���            B  �  �  O         ����   J K          � '�� y     �  �x  $!   ��  �       ���            C  �  �  O         ����   M O          � -�� z     �  z  l3   ��  �       ���            D  �  �  O         ����   S T          � 3�� {       �{  �E   ��  �       ���            E  �  �  O         ����   W Y          � 9� |     >  �|  �W   ��  �       ���            F  �  �  O         ����   [ ]          � ?
� }     m  T~  Dj   ��  �       ���            G  �  �  O         ����   J L          � ?� �     m  ��  ��   ��  �
       ���            "L  �  �  P         ����   N O          � E� �     �  F�  ԫ   ��  �       ���            !M  �  �  P         ����   R S          � K!� �     �  ̍  (�   ��  �       ���             N  �  �  P         ����   X Y          � Q)� �       R�  |�   ��  �       ���            O  �  �  P         ����   \ ^          � W1� �     I  ؐ  ��   ��  �       ���            P  �  �  P         ����   a b          ]9� �     �  ^�  $   ��  �       ���            Q  �  �  P         ����   P Q          ]@� �     �  ��  �[	   ��  �
       ��{            .L  �  �           ����   T U          cH� �     4  ^�  �t	   ��  �       ��{            -M  �  �           ����   X Y          iP� �     s  �  �	   ��  �       ��{            ,N  �  �           ����   ^ `          oX� �     �  ��  ��	   ��  �       ��{            +O  �  �           ����   c d          $u`� �     �  J�  V�	   ��  �       ��{            *P  �  �           ����   h i          *{h� �     0  �  ��	   ��  �       ��{            )Q  �  �           ����   T U          ,�n�     (  :�  �c   ��  �
       ��|            ;V  �  �           ����   X Y          2�v�     p  ��  �   ��  �       ��|            :W  �  �           ����   \ ^          8�~�     �  ��  ��   ��  �       ��|            9X  �  �           ����   c d          >���        ��   �   ��  �       ��|            8Y  �  �           ����   h i          D���     H  B�   �   ��  �       ��|            7Z  �  �           ����   m o          J�� �     �  �  @�   ��  �       ��|            6[  �  �           ����   9 :          | � Ff       �  h=  �(      �
     �   �            � .  �  �  X         ����   < =          � � Mj       �  X>  1       �     �   �            � /  �  �  X         ����   ? @          � � Tn       �  H?  �9   ��  �     �   �            � 0  �  �  X         ����   C D          � � [r       �  8@  �A   ��  �     �   �            � 1  �  �  X         ����   F H          � � bv       �  (A  hJ   ��  �     �   �            � 2  �  �  X         ����   J K          � � iz       �  B  �R   ��  �     �   �            � 3  �  �  X         ����   = >          � � ou       z  �J  ��   ��  �
     �   �           	 � 8  �  �  Y         ����   @ A          � � vy       �  �K  4�   ��  �     �   �           	 � 9  �  �  Y         ����   C D          � � }}       �  �L  �    ��  �     �   �           	 � :  �  �  Y         ����   H I          � � ��       �  �M  L   ��  �     �   �           	 � ;  �  �  Y         ����   K M          � � ��       �  �N  �   ��  �     �   �           	 � <  �  �  Y         ����   O Q          � � ��         
P  d    ��  �     �   �           	 � =  �  �  Y         ����   ? A          � � ��       �	  �Y  "�   ��  �
     �   �           
 8  �  �  Z         ����   C D          � � ��       �	  �Z  �   ��  �     �   �           
 9  �  �  Z         ����   F G          � � ��       
  �[  ��   ��  �     �   �           
 :  �  �  Z         ����   K L          � � ��       ?
  *]  �    ��  �     �   �           
 ;  �  �  Z         ����   O P          � � ��       `
  V^  �   ��  �     �   �           
  <  �  �  Z         ����   S T          � � ��       �
  �_  �   ��  �     �   �           
 � =  �  �  Z         ����   D E          � �� n     �  j  ��   ��  �
     �   �            B  �  �  [         ����   G H          � �� o     �  Xk      ��  �     �   �            C  �  �  [         ����   J L          � �� p     
  �l  �   ��  �     �   �            D  �  �  [         ����   P Q          � �� q     2  �m  '   ��  �     �   �            
E  �  �  [         ����   T U          � �� r     Z  6o  �6   ��  �     �   �            	F  �  �  [         ����   X Z          �  �� s     �  �p   F   ��  �     �   �            G  �  �  [         ����   H I          � !�� x       �{  �K   ��  �
     �   �            B  �  �  \         ����   K M          � '�� y     M  d}  ^   ��  �     �   �            C  �  �  \         ����   O P          � -�� z     |  �~  \p   ��  �     �   �            D  �  �  \         ����   T V          � 3� {     �  4�  ��   ��  �     �   �            E  �  �  \         ����   Y Z          � 9� |     �  ��  �   ��  �     �   �            F  �  �  \         ����   ] _          � ?� }     	  �  4�   ��  �     �   �            G  �  �  \         ����   L M          � ?� �       p�   �   ��  �
     �   �            "L  �  �  ]         ����   O Q          � E%� �     L  ��  t�   ��  �     �   �            !M  �  �  ]         ����   S U          � K-� �     �  |�  �   ��  �     �   �             N  �  �  ]         ����   Y [          � Q5� �     �  �     ��  �     �   �            O  �  �  ]         ����   ^ _          � W=� �     �  ��  p-   ��  �     �   �            P  �  �  ]         ����   b d          ]E� �     (  �  �B   ��  �     �   �            Q  �  �  ]         ����   Q R          ]L� �     �  j�  6�	   ��  �
     �   �            .L  �  �           ����   U V          cT� �     �  �  Һ	   ��  �     �   �            -M  �  �           ����   Y [          i\� �     '  ��  n�	   ��  �     �   �            ,N  �  �           ����   ` a          od� �     f  V�  
�	   ��  �     �   �            +O  �  �           ����   d f          $ul� �     �  ��  �
   ��  �     �   �            *P  �  �           ����   i k          *{t� �     �  ��  B
   ��  �     �   �            )Q  �  �           ����   T U          ,�z�     �  �  ��   ��  �
     �   �            ;V  �  �           ����   X Y          2���     0  ��  ��   ��  �     �   �            :W  �  �           ����   \ ^          8���     x  n�  ��   ��  �     �   �            9X  �  �           ����   c d          >���     �  0�      ��  �     �   �            8Y  �  �           ����   h i          D���       ��      ��  �     �   �            7Z  �  �           ����   m o          J�� �     P  ��  @;   ��  �     �   �            6[  �  �            ��� ��     
                     ��     �     �
  !  �� ���        ������  ����������������        ��� ��     
                     ��     �     �
  "  �� ���        ������  ����������������        ��� ��     
                     ��     �     �
  #  �� ���        ������  ����������������        ��� ��                          ��     �     �
  $  �� ���        ������  ����������������        ��� ��                          ��     �     �
  %  �� ���        ������  ����������������        ��� ��                          ��     �     �
  &  �� ���        ������  ����������������        ��� ��     (                     ��     �     �
  '  �� ���        ������  ����������������        ��� ��     (                     ��     �     �
  (  �� ���        ������  ����������������        ��� ��     (                     ��     �     �
  )  �� ���        ������  ����������������        ��� ��   m 2                     ��     �     �
    �� ���        ������  ����������������        ��� ��  
                         �  �� �     �
    �� ���        ������  ����������������        ��� �� ( 
                         �   � �     �
    �� ���        ������  ����������������        ��� �� < 
                         �  @B �     �
    �� ���        ������  ����������������        ��� �� d   �                         �     �     �
    ! ���        ������  ����������������        ��� �� d   �                         �     �     �
     ���        ������  ����������������        ��� �� d   �                         �     �     �
      ���        ������  ����������������        ��� ��	 d   �                         �     �     �
    " ���        ������  ����������������        ��� ��                            ��     �     �
    �� ���        ������  ����������������        ��� ��                            ��     �     �
  *  �� ���        ������  ����������������        ��� ��                            ��     �     �
  +  �� ���        ������  ����������������        ��� ��                         ��     �     �
    �� ���        ������  ����������������        ��� ��                         ��     �     �
  ,  �� ���        ������  ����������������        ��� ��                         ��     �     �
  -  �� ���        ������  ����������������        ��� ��                         ��     �     �
    �� ���        ������  ����������������        ��� ��                         ��     �     �
  ,  �� ���        ������  ����������������        ��� ��                         ��     �     �
  -  �� ���        ������  ����������������        �� �  d d x   

-                    �  '  �     �
     ��y ���        ������  ����������������        �� �    x   

-                    @  �8 �     �
      ��z ���        ������  ����������������        �����                                 �   �  �     �
  !   �� ���        ������  ����������������       ��  � ��    %                                        �
      ��{ ���        ������  ����������������       ��  � ��    &                                        �
      ��{ ���        ������  ����������������       ��  � ��    '                                        �
      ��{ ���        ������  ����������������       ��  � ��    (                                        �
      ��{ ���        ������  ����������������       ��  � ��    )                                        �
      ��{ ���        ������  ����������������       �� � ��    �F   �F                                  �
      ��{ ���        ������  ����������������       �� � ��    �F   �F                                  �
      ��{ ���        ������  ����������������       �� � ��    �F   �F                                  �
      ��{ ���        ������  ����������������       �� � ��    �F   �F                                  �
      ��{ ���        ������  ����������������       �� � ��    �F   �F                                  �
      ��{ ���        ������  ����������������       �� � ��� ��F   �F                                  �
      ��{ ���        %   ��  ����������������       �� � �����F   �F                                  �
      ��{ ���        %   ��  ����������������       �� � �����F   �F                                  �
      ��{ ���        %   ��  ����������������       �� � ���T�F   �F                                  �
      ��{ ���        %   ��  ����������������       �� � ��`	�F   �F                                  �
      ��{ ���        %   ��  ����������������        ��p ��  3                        �����  �        �
     ��, ���        ������  ����������������        ��p ��  9                        �����  �        �
     ��, ���        ������  ����������������        ��p ��  ?                        �����  �        �
     ��, ���        ������  ����������������        ��p ��  ,                        �����  �        �
     ��, ���        ������  ����������������        ��p ��  j                        �����  �        �
     ��, ���        ������  ����������������        ����� ��                               �  '  �     �
  "   �� ��x        ������  ����������������        ����� ��                               �   N  �     �
  "   �� ��}        ������  ����������������        ����� ��                               @  ��  �     �
  "   �� ��Q        ������  ����������������        ����� ��                               �.  ��  �     �
  "   �� ��L        ������  ����������������        ����� ��                               �>  �8 �     �
  "   �� ��r        ������  ����������������        � g                 �$��n     ������  %�       �
      ��) ��U        ����   ����������������        � g                 �L��}     ����h�  �       �
      ��) ��U        ����   ����������������          ��I��2    � <��         ȇ  �l      d 
     `   �     Y#V#    �   �  �  �             ����x2    � B��       7  N�  D�      d      `   �     Y#V#    �   �  �  �             ���A\�2    � H �       m  Ԋ  ��      d      `   �     Y#V$    �   �  �  �             ����`2    � N�       �  Z�  �      d      `   �     Y#V$    �   �  �  �             ��c�@�2    � T�       �  ��  @�      d      `   �     Y#V"    �   �  �  �             ���N�M2    Z�         f�  ��      d      `   �     Y#V"    �   �  �  �           ��p ��  3                        �����  �  �    �
     ��, ���        ������  ����������������        ��p ��  9                        �����  �  �    �
     ��, ���        ������  ����������������        ��p ��  ?                        �����  �  �    �
     ��, ���        ������  ����������������        ��p ��  ,                        �����  �  �    �
     ��, ���        ������  ����������������        ��p ��  j                        �����  �  �    �
     ��, ���        ������  ����������������          ���w�o2    �Z� �       @   }   Y                 �     �m�    �    �  �  �             ��g�t2    �`� �       o  h~  Hk                 �     �m�    � 	   �  �  �             ����)�2    �f� �       �  �  �}                 �     �m�    � �����  �  �             ���C�W2    w� �       S  (�  0�                 �    TX�    
   �  �  �             ��1�Y 2    #}� �       �  ��  �                 �    TX�    		   �  �  �             ����(�2    +�� �       �  4�  �                 �    TX�    �����  �  �             ��f�Q2    J�         ֦  ��	   ��            �    :��    �    �  �  �             ����U	2    R�      E  z�  &�	   ��            �    :��    �    �  �  �             ����@	
2    Z�
      �  �  ��	   ��            �    :��    � �����  �  �             ��=��l	2    x�2&      h  
�  ��   ��            �    �Z       �  �  �             ����l	E
2    ��8,      �  ̿  ��   ��            �    �Z       �  �  �             ����	u
f2    ��>2      �  ��  �   ��            �    �Z    �����  �  �             ����	�
2    ��RFt     �$  ��  C   ��            �   ���       �  �  �            ����	�
t2    ��XLu     �$  ��  �b   ��            �   ���       �  �  �            ���	�
��2    ��^Rv     #%  ��  Ă   ��            �   ���     �����  �  �            ����	�
�2    �qe~     b+  �  H�   ��            �   ���       �  �  �            ���	�
��2    �wk     �+  �  $   ��            �   ���       �  �  �            ���
�$2    �!}q�     ,   �   :   ��            �   ���    �����  �  �            ���	�
��2    G���     3  � ��   ��               ���    &   �  �  �            ���
��'2    O���     y3  �    ��               ���    '   �  �  �            ���Hd�2    (W���     �3   &C   ��               ���    �����  �  �            ���
G2    Jt���     �;  * �I   ��            '   ���    *&   �  �  �            ���-L�2    S|���     <  P, @v   ��            '   ���    )'   �  �  �            ��)��F2    \����     �<  �. Ȣ   ��            '   ���    (�����  �  �            ���<e�2    }����     E  �H �   ��            (   ���    0   �  �  �            ���m�2    �����     �E  @K @,   ��            (   ���    1   �  �  �            ��lk�2    �����     F  �M x]   ��            (   ���    �����  �  �            ���S��2    ��."�     �;  * �I   ��  �
     �    �   ���    0   �  �  �            ����]2    ��5)�     <  P, @v   ��  �
     �    �   ���    1   �  �  �            ������2    ��<0�     �<  �. Ȣ   ��  �
     �    �   ���    �����  �  �            ��k_(�2    ��."�     E  �H �   ��  �
     �    �   ���    0   �  �  �            ����2    ��5)�     �E  @K @,   ��  �
     �    �   ���    1   �  �  �            ��p��2    ��<0�     F  �M x]   ��  �
     �    �   ���    �����  �  �            ��W�z
2    �i� �       `  �}  0e       #      !   �    �}Y    � :   �  �  �             �����2    �o� �       �  X  xw       #      !   �    �}Y    � ;   �  �  �             ���_k2    u� �       �  ��  ��       #      !   �    �}Y    � �����  �  �             ��F�$�2    *�� �       o  �  P�       $      "   �    P�b    
:   �  �  �             �����Q2    2�� �       �  ��  �       $      "   �    P�b    	;   �  �  �             ����	82    :�� �       �  $�  �'       $      "   �    P�b    �����  �  �             ��:���2    Y�       *  Ƨ  ��	   ��  %      #   �    66�    � D   �  �  �             ����	S!2    a�      i  j�  6�	   ��  %      #   �    66�    � E   �  �  �             ���	�
�2    i�
      �  �  �
   ��  %      #   �    66�    � �����  �  �             ��M	
�W2    ��2&      �  ��  ��   ��  &      $   �    ��    D   �  �  �             ��#
 2    ��8,      �  ��  �   ��  &      $   �    ��    E   �  �  �             ��A>��2    ��>2        ~�  �'   ��  &      $   �    ��    �����  �  �             ��n
U?32    ��RFt     �$  ��  �R   ��  '      %   �   ���    N   �  �  �            ��^Z��2    �XLu      %  ��  �r   ��  '      %   �   ���    O   �  �  �            ������	2    �^Rv     R%  t�  ��   ��  '      %   �   ���     �����  �  �            ����	2    �"qe~     �+  ��  (   ��  (      &   �   ���    N   �  �  �            ������	2    �)wk     �+  ��  '   ��  (      &   �   ���    O   �  �  �            ��L�	 2    0}q�     F,  ��  �J   ��  (      &   �   ���    �����  �  �            ���
�
2    %V���     B3  � �   ��  )      '      ���    X   �  �  �            ��N�	�
2    .^���     �3  � �,   ��  )      '      ���    Y   �  �  �            �����
2    7f���     4  � �T   ��  )      '      ���    �����  �  �            ��?u�		2    Y����     �;  + x\   ��  *      (   )   ���    *X   �  �  �            �����
2    b����     @<  @-  �   ��  *      (   )   ���    )Y   �  �  �            ��<��Z2    k����     �<  z/ ��   ��  *      (   )   ���    (�����  �  �            �����
2    �����     DE  �I �   ��  +      )   *   ���    b   �  �  �            ��x�$2    �����     �E  0L �?   ��  +      )   *   ���    c   �  �  �            ������2    �����     @F  �N (q   ��  +      )   *   ���    �����  �  �            ���?�2    ��."�     �;  + x\   ��  �
     �   �   ���    b   �  �  �            ��x?C"2    �5)�     @<  @-  �   ��  �
     �   �   ���    c   �  �  �            �����2    �<0�     �<  z/ ��   ��  �
     �   �   ���    �����  �  �            ���I�2    ��."�     DE  �I �   ��  �
     �   �   ���    b   �  �  �            ���KJ)2    �5)�     �E  0L �?   ��  �
     �   �   ���    c   �  �  �            �����2    �<0�     @F  �N (q   ��  �
     �   �   ���    �����  �  �            ��pp2    �� ��       I  <}  \       7      5   �    �V#    � l   �  �  �             ������2    �� ��       x  �~  Tn       7      5   �    �V#    � m   �  �  �             ���F�F2    �� ��       �  �  ��       7      5   �    �V#    � �����  �  �             ��4�4�2    �� ��       V  d�  x�       8      6   �    ��H    
l   �  �  �             ���z�z2    ���       �  �  �       8      6   �    ��H    	m   �  �  �             ���L�L2    ���       �  p�          8      6   �    ��H    �����  �  �             ����2            �  �	   ��  9      7   �    <|�    � v   �  �  �             ����2    

      N  ��  ��	   ��  9      7   �    <|�    � w   �  �  �             ���n	�n	2          �  Z�  F�	   ��  9      7   �    <|�    � �����  �  �             ������2    8:8.      q  F�  `�   ��  :      8   �    ׂ�    v   �  �  �             ����	��	2    @@@4      �  �  �    ��  :      8   �    ׂ�    w   �  �  �             ���	�
�	�
2    HFH:        ��  �   ��  :      8   �    ׂ�    �����  �  �             ����	��	2    fZfNt     �$   �   G   ��  ;      9   �   ���    �   �  �  �            ���	�
�	�
2    n`nTu     �$  ��  �f   ��  ;      9   �   ���    �   �  �  �            ���
��
�2    vfvZv     *%  ��  ��   ��  ;      9   �   ���     �����  �  �            ���	�
�	�
2    �y�m~     n+  @�  ��   ��  <      :   �   ���    �   �  �  �            ���
��
�2    ��s     �+  >�  \   ��  <      :   �   ���    �   �  �  �            ���&�&2    ���y�     &,  <�  8>   ��  <      :   �   ���    �����  �  �            ���
�
2    �����      3   r�   ��  =      ;      ���    �   �  �  �            ����2    �����     �3  " �   ��  =      ;      ���    �   �  �  �            ��@�@�2    �����     �3  > �G   ��  =      ;      ���    �����  �  �            ��FF2    �����     �;  R* hN   ��  >      <   +   ���    *�   �  �  �            ��$x$x2    ���     <  �, �z   ��  >      <   +   ���    )�   �  �  �            ����2    ���     �<  �. x�   ��  >      <   +   ���    (�����  �  �            ��:�:�2    0�0��     E  $I ��   ��  ?      =   ,   ���    �   �  �  �            ��j�j�2    9�9��     �E  |K ,1   ��  ?      =   ,   ���    �   �  �  �            �� � �2    B�B��     F  �M db   ��  ?      =   ,   ���    �����  �  �            ��^^2    �6�*�     �;  R* hN   ��  �
     �   �   ���    �   �  �  �            ������2    �=�1�     <  �, �z   ��  �
     �   �   ���    �   �  �  �            ��2    �D�8�     �<  �. x�   ��  �
     �   �   ���    �����  �  �            ��ff2    �6�*�     E  $I ��   ��  �
     �   �   ���    �   �  �  �            ������2    �=�1�     �E  |K ,1   ��  �
     �   �   ���    �   �  �  �            ��2    �D�8�     F  �M db   ��  �
     �   �   ���    �����  �  �            ���o�w2    �d� �       Q  �}  $b       M      J   �    C�!    � �   �  �  �             ��tg�2    �j� �           lt       M      J   �    C�!    � �   �  �  �             ��)���2    �p� �       �  ��  ��       M      J   �    C�!    � �����  �  �             ���W�C2    %�� �       n  ܑ  �       N      K   �    �s�!    
�   �  �  �             ��Y 1�2    -�� �       �  b�  \       N      K   �    �s�!    	�   �  �  �             ��(���2    5�� �       �  �  �$       N      K   �    �s�!    �����  �  �             ���Qf2    T�       !  ��  �	       O      L   �    ��H!    � �   �  �  �             ��U	��2    \�      `  .�  ��	       O      L   �    ��H!    � �   �  �  �             ��@	
��2    d�
      �  Ҫ  N
       O      L   �    ��H!    � �����  �  �             ���l	=�2    ��2&      �  ��  ��       P      M   �    ���!    �   �  �  �             ��l	E
��2    ��8,      �  ��          P      M   �    ���!    �   �  �  �             ��u
f��	2    ��>2        B�   $       P      M   �    ���!    �����  �  �             ���	�
�2    ��RFt     �$  x�  �N       Q      N   �   ���!    �   �  �  �            ���
t��	2    � XLu     �$  X�  �n       Q      N   �   ���!    �   �  �  �            �����	�
2    �^Rv     H%  8�  ��       Q      N   �   ���!     �����  �  �            ���
���	2    �qe~     |+  ��  ��       R      O   �   �ؓ!    �   �  �  �            �����	�
2    �$wk     �+  ��  �"       R      O   �   �ؓ!    �   �  �  �            ��$�
�2    �+}q�     2,  ��  �F       R      O   �   �ؓ!    �����  �  �            �����	�
2     Q���     /3  ~ Z        S      P      ���!    �   �  �  �            ���'�
�2    )Y���     �3  � n(       S      P      ���!    �   �  �  �            ��d��H2    2a���     �3  � �P       S      P      ���!    �����  �  �            ��G�
2    T~���     �;  �* �W       T      Q   -   ���!    *�   �  �  �            ��L��-2    ]����     4<  - P�       T      Q   -   ���!    )�   �  �  �            ���F)�2    f����     �<  >/ ذ       T      Q   -   ���!    (�����  �  �            ��e��<2    �����     7E  �I �	       U      R   .   ���!    �   �  �  �            ����m2    �����     �E  �K ;       U      R   .   ���!    �   �  �  �            ��k�l2    �����     3F  LN <l       U      R   .   ���!    �����  �  �            �����S2    ��."�     �;  �* �W       �
     �   �   ���!    �   �  �  �            ���]�2    �5)�     4<  - P�       �
     �   �   ���!    �   �  �  �            ������2    �	<0�     �<  >/ ذ       �
     �   �   ���!    �����  �  �            �����\2    ��."�     7E  �I �	       �
        �   ���!    �   �  �  �            ���g�2    �5)�     �E  �K ;       �
        �   ���!    �   �  �  �            ����� 2    �	<0�     3F  LN <l       �
        �   ���!    �����  �  �            ��z
W�2    � B��       9  �|  �U       c      _   �    Cc!    � �   �  �  �             �����2    � H��       h  ,~  <h       c      _   �    Cc!    � �   �  �  �             ��k�_2    � N��       �  �  �z       c      _   �    Cc!    � �����  �  �             ��$�F�2    ` �       E  �  ��      d      `   �     Y#V!    
�   �  �  �             ���Q��2    f(�       {  r�  <      d      `   �     Y#V!    	�   �  �  �             ��8��	2    l0�       �  ��  �      d      `   �     Y#V!    �����  �  �             ����:�2    -~O      �  ��  �	       e      a   �    �y !    � �   �  �  �             ��S!��	2    3�W      <  >�  ��	       e      a   �    �y !    � �   �  �  �             ����	�
2    9�_      {  �  >�	       e      a   �    �y !    � �����  �  �             ���WM	
2    M�},      ^  ν  ��       f      b   �    ��!    �   �  �  �             �� #
2    S��2      �  ��   �       f      b   �    ��!    �   �  �  �             ����A>2    Y��8      �  R�          f      b   �    ��!    �����  �  �             ��?3n
U2    m��Lt     {$  ��  ?       g      c   �   ���!    �   �  �  �            ����^Z2    s��Ru     �$  h�  �^       g      c   �   ���!    �   �  �  �            ����	��2    y��Xv     %  H�  �~       g      c   �   ���!     �����  �  �            ��	��2    ���k~     X+  ��  �       h      d   �   ��X!    �   �  �  �            ����	��2    ���q     �+  ��  �       h      d   �   ��X!    �   �  �  �            ���	 L2    ��w�     ,  ��  �5       h      d   �   ��X!    �����  �  �            ���
�
2    ���     	3  � ��       i      e      ���!    �   �  �  �            ���	�
N2    �#$��     p3  � �       i      e      ���!    �   �  �  �            ���
��2    �*-��     �3  � �>       i      e      ���!    �����  �  �            ���		?u2    �PO��     �;  �) E       j      f   /   ���!    *�   �  �  �            ���
��2    �XX��     <  , �q       j      f   /   ���!    )�   �  �  �            ���Z<�2    �`a��     v<  N. �       j      f   /   ���!    (�����  �  �            ���
��2    ~���     E  �H �       k      g   0   ���!    �   �  �  �            ���$x2    ����     �E  K T'       k      g   0   ���!    �   �  �  �            ������2    ����     F  \M �X       k      g   0   ���!    �����  �  �            ����?2    S��(�     �;  �) E       �
       �   ���!    �   �  �  �            ��C"x?2    Z��/�     <  , �q       �
       �   ���!    �   �  �  �            �����2    a��6�     v<  N. �       �
       �   ���!    �����  �  �            ����I2    S��(�     E  �H �       �
       �   ���!    �   �  �  �            ��J)�K2    Z��/�     �E  K T'       �
       �   ���!    �   �  �  �            �����2    a��6�     F  \M �X       �
       �   ���!    �����  �  �             0�0�
2    �� ��       Q  x}  _       }      w   �    ���    �   �  �  �              �:�:
2    �� ��       �  �~  `q       }      w   �    ���    �   �  �  �              G�G�
2    �� ��       �  H�  ��       }      w   �    ���    � �����  �  �              ����
2    �� ��       f  ��  ��       ~      x   �    ���    
  �  �  �              oo
2    ���       �  &�         ~      x   �    ���    	  �  �  �              $�$�
2    ���       �  ��  h!       ~      x   �    ���    �����  �  �              �b�b
2            N�  ��	             y   �    ���    �   �  �  �              NN
2    
      W  �  .�	             y   �    ���    �   �  �  �              ��
2          �  ��  ��	             y   �    ���    � �����  �  �              �X�X
2    6:8.      {  ��   �       �      z   �    ���      �  �  �              3	3	
2    >@@4      �  D�  @       �      z   �    ���      �  �  �              	
	

2    FFH:        �  `        �      z   �    ���    �����  �  �              mT	mT	
2    dZfNt     �$  <�  �J       �      {   �   ���      �  �  �             /	+
/	+

2    l`nTu     �$  �  �j       �      {   �   ���      �  �  �             2
J2
J
2    tfvZv     4%  ��  ��       �      {   �   ���     �����  �  �             Y	e
Y	e

2    �y�m~     y+  |�  ��       �      |   �   ���      �  �  �             0
U0
U
2    ��s     �+  z�  �       �      |   �   ���      �  �  �             O�O�
2    ���y�     1,  x�  pB       �      |   �   ���    �����  �  �             _
�_
�
2    �����     +3  B ��       �      }      ���       �  �  �             N�N�
2    �����     �3  ^ �#       �      }      ���    !  �  �  �             ����
2    �����     �3  z L       �      }      ���    �����  �  �             h�h�
2    �����     �;  �* S       �      ~   1   ���    *   �  �  �             o�o�
2    ���     (<  �, �       �      ~   1   ���    )!  �  �  �             �W�W
2    ���     �<  / (�       �      ~   1   ���    (�����  �  �             ����
2    .�0��     +E  `I �       �         2   ���    *  �  �  �             ��
2    7�9��     �E  �K 6       �         2   ���    +  �  �  �             #�#�
2    @�B��     'F  N Pg       �         2   ���    �����  �  �             o'o'
2    �6�*�     �;  �* S       �
       �   ���    *  �  �  �             ����
2    �=�1�     (<  �, �       �
       �   ���    +  �  �  �             ����
2    �D�8�     �<  / (�       �
       �   ���    �����  �  �             y0y0
2    �6�*�     +E  `I �       �
       �   ���    *  �  �  �             ����
2    �=�1�     �E  �K 6       �
       �   ���    +  �  �  �             ��
2    �D�8�     'F  N Pg       �
       �   ���    �����  �  �             �z
2    k�� �       _  �}  0e       �      �       ���    �    �  �  �             �9�2    q�� �       �  X  xw       �      �       ���    � 	   �  �  �             Ck2    w�� �       �  ��  ��       �      �       ���    � �����  �  �             ��$�2    ��� �       o  �  P�       �      �   	   ioe    
   �  �  �             �E�Q2    ��� �       �  ��  �       �      �   	   ioe    		   �  �  �             W.	82    ��� �       �  $�  �'       �      �   	   ioe    �����  �  �             ����2    �%       *  Ƨ  ��	       �      �   
   ��    �    �  �  �             �n	S!2    �-      i  j�  6�	       �      �   
   ��    �    �  �  �             �	x
�2    �5
      �  �  �
       �      �   
   ��    � �����  �  �             ��	�W2    �T2&      �  ��  ��       �      �      :��       �  �  �             �	�
 2    �\8,      �  ��  �       �      �      :��       �  �  �             �
���2    �d>2        ~�  �'       �      �      :��    �����  �  �             �	�
?32    �RFt     �$  ��  �R       �      �   �   ���       �  �  �             �
���2    �XLu      %  ��  �r       �      �   �   ���       �  �  �             @��	2    �^Rv     R%  t�  ��       �      �   �   ���     �����  �  �             0	2    9�qe~     �+  ��  (       �      �   �   ���       �  �  �             I��	2    A�wk     �+  ��  '       �      �   �   ���       �  �  �             g��	 2    I�}q�     F,  ��  �J       �      �   �   ���    �����  �  �             G��
2    e����     B3  � �       �      �      ���    &   �  �  �             a��	�
2    m����     �3  � �,       �      �      ���    '   �  �  �             �_�
2    u����     4  � �T       �      �      ���    �����  �  �             ���		2    �!���     �;  + x\       �      �   3   ���    *&   �  �  �             �9�
2    �*���     @<  @-  �       �      �   3   ���    )'   �  �  �             a�Z2    �3���     �<  z/ ��       �      �   3   ���    (�����  �  �             �R�
2    �V���     DE  �I �       �      �   4   ���    0   �  �  �             >��$2    �_���     �E  0L �?       �      �   4   ���    1   �  �  �             ���2    �h���     @F  �N (q       �      �   4   ���    �����  �  �             �m�2    	�."�     �;  + x\       �
       �   ���    0   �  �  �             {ZC"2    �5)�     @<  @-  �       �
       �   ���    1   �  �  �             ���2    �<0�     �<  z/ ��       �
       �   ���    �����  �  �             �u�2    	�."�     DE  �I �       �
       �   ���    0   �  �  �             �dJ)2    �5)�     �E  0L �?       �
       �   ���    1   �  �  �             ���2    �<0�     @F  �N (q       �
       �   ���    �����  �  �         ����   c e          y� � ~       �  86  ��             ��            � 4  �  �  �          ����   n q          �� � �       �  86  ��             ��            � 5  �  �  �          ����   ~ �          �� � �       �  86  ��             ��            � �����  �  �          ����   j m          �� � �       |  �J  p�            	  ��	           	 � >  �  �  �          ����   w z          �� � �       �  �K  ��            	  ��	           	 � ?  �  �  �          ����   � �          �� �       �  �L  �            	  ��	           	 � �����  �  �          ����   p r          �� �       �	  nZ  ��   ��       
  ��           
 � >  �  �  �         ����   } �          �$� �       
  �[  ��   ��       
  ��           
 � ?  �  �  �         ����   � �          �*� �       4
  �\  ��   ��       
  ��           
 � �����  �  �         ����   x z          �=� � t     �  �k  x
   ��          ���            H  �  �  �         ����   � �          �C� � u       �l  �   ��          ���            I  �  �  �         ����   � �          �I� � v     :  n  h)   ��          ���            �����  �  �         ����   ~           '[� � ~     h  ,~  <h   ��  !       ���            H  �  �  y         ����   � �          /a� �      �  �  �z   ��  !       ���            I  �  �  y         ����   � �          7g� � �     �  ��  ̌   ��  !       ���            �����  �  y         ����   � �          Vx� � �       T�  �    ��  "       ��'            R  �  �  �         ����   � �          ^~� � �     �  ړ  �   ��  "       ��'            S  �  �  �         ����   � �          f�� � �     �  `�  @+   ��  "       ��'            �����  �  �         ����   � �          �� �     3  �  �	   ��  #       ��5            (R  �  �  �         ����   � �          ���     r  ��  ��	   ��  #       ��5            'S  �  �  �         ����   � �          ��
�     �  J�  V	
   ��  #       ��5            &�����  �  �         ����   � �          ��2&�     �  6�  `�   ��  $       ��6            5\  �  �  �         ����   � �          ��8,�     �  ��  �   ��  $       ��6            4]  �  �  �         ����   � �          ��>2�     (  ��  �+   ��  $       ��6            3�����  �  �         ����  ` c          3� n b       �  D4  d�   ��  �       ��            � 4  �  �  �          ����  l n          3� n b       �  D4  d�   ��  �       ��            � 5  �  �  �          ����  { ~          3� n b       �  D4  d�   ��  �       ��            � �����  �  �          ����  g h          �� � �       J  �H  ��   ��  �     	  ��           	 � >  �  �  �          ����  s u          �� � �       e  �I  t�   ��  �     	  ��           	 � ?  �  �  �          ����  � �          �� �       �   K   �   ��  �     	  ��           	 � �����  �  �          ����  o p          �� �       �	  zX  >�   ��  �     
  ��           
 � >  �  �  �         ����  | }          �$� �       �	  �Y  "�   ��  �     
  ��           
 � ?  �  �  �         ����  � �          �*� �       �	  �Z  �   ��  �     
  ��           
 � �����  �  �         ����  t v          �=� � t     �  �i  �   ��  �       ���            H  �  �  �         ����  � �          �C� � u     �  �j  �   ��  �       ���            I  �  �  �         ����  � �          �I� � v     �  *l  �   ��  �       ���            �����  �  �         ����  | ~          [� � ~     '  8|  �N   ��  �       ���            H  �  �  {         ����  � �          a� �      V  �}   a   ��  �       ���            I  �  �  {         ����  � �          "g� � �     �    hs   ��  �       ���            �����  �  {         ����  � �          Ax� � �     9  `�  @�   ��  �       ��,            R  �  �  �         ����  � �          I~� � �     p  �  ��   ��  �       ��,            S  �  �  �         ����  � �          Q�� � �     �  l�  �   ��  �       ��,            �����  �  �         ����  � �          p� �     �  �  Һ	   ��  �       ��A            (R  �  �  �         ����  � �          x��     '  ��  n�	   ��  �       ��A            'S  �  �  �         ����  � �          ��
�     f  V�  
�	   ��  �       ��A            &�����  �  �         ����  � �          ��2&�     H  B�   �   ��  �       ��B            5\  �  �  �         ����  � �          ��8,�     �  �  @�   ��  �       ��B            4]  �  �  �         ����  � �          ��>2�     �  ��  `   ��  �       ��B            3�����  �  �         ����  c e          q� � ~       E  p:  �   ��  �       ��A            � 4  �  �           ����  n q          x� � �       [  `;  `   ��  �       ��A            � 5  �  �           ����  ~ �          � � �       q  P<  �   ��  �       ��A            � �����  �           ����  h j          �� � �       @  �H   �   ��  �     	  ��B           	 � >  �  �           ����  u w          �� � �       [  �I  ��   ��  �     	  ��B           	 � ?  �  �           ����  � �          �� �       v  �J  �   ��  �     	  ��B           	 � �����  �           ����  p r          �� �       �	  X  ��   ��  �     
  ��           
 � >  �  �  �         ����  } �          �$� �       �	  BY  ��   ��  �     
  ��           
 � ?  �  �  �         ����  � �          �*� �       �	  nZ  ��   ��  �     
  ��           
 � �����  �  �         ����  v x          �=� � t     �  2i  X�   ��  �       ���            H  �  �  �         ����  � �          �C� � u     �  |j  ��   ��  �       ���            I  �  �  �         ����  � �          �I� � v     �  �k  H   ��  �       ���            �����  �  �         ����  ~           [� � ~       �{  �I   ��  �       ���            H  �  �  z         ����  � �          'a� �      I  <}  \   ��  �       ���            I  �  �  z         ����  � �          /g� � �     x  �~  Tn   ��  �       ���            �����  �  z         ����  � �          Nx� � �     +  ��  ��   ��  �       ��2            R  �  �  �         ����  � �          V~� � �     b  ��  �   ��  �       ��2            S  �  �  �         ����  � �          ^�� � �     �  �  p
   ��  �       ��2            �����  �  �         ����  � �          }� �     �  ��  ��	   ��  �       ��M            (R  �  �  �         ����  � �          ���       N�  ��	   ��  �       ��M            'S  �  �  �         ����  � �          ��
�     W  �  .�	   ��  �       ��M            &�����  �  �         ����  � �          ��2&�     8  ޼  ��   ��  �       ��N            5\  �  �  �         ����  � �          ��8,�     �  ��   �   ��  �       ��N            4]  �  �  �         ����  � �          ��>2�     �  b�      ��  �       ��N            3�����  �  �         ����  ` c          _� � ~       �  xA  8M   ��  ]       ��T            � 4  �  �            ����  l n          f� � �       �  hB  �U   ��  ]       ��T            � 5  �  �            ����  { ~          m� � �         XC  ^   ��  ]       ��T            � �����  �            ����  g h          �� � �       �  �O  P   ��  ^     	  ��U           	 � >  �  �  !         ����  s u          �� � �         �P  �%   ��  ^     	  ��U           	 � ?  �  �  !         ����  � �          �� �       *  �Q  h0   ��  ^     	  ��U           	 � �����  �  !         ����  o p          �� �       v
  _  J   ��  _     
  ��           
 � >  �  �  �         ����  | }          �$� �       �
  J`  .#   ��  _     
  ��           
 � ?  �  �  �         ����  � �          �*� �       �
  va  0   ��  _     
  ��           
 � �����  �  �         ����  t v          �=� � t     z  :p  �B   ��  `       ���            H  �  �  �         ����  � �          �C� � u     �  �q  0R   ��  `       ���            I  �  �  �         ����  � �          �I� � v     �  �r  �a   ��  `       ���            �����  �  �         ����  | ~          [� � ~       ܂  ,�   ��  a       ���            H  �  �  |         ����  � �          a� �      3  D�  t�   ��  a       ���            I  �  �  |         ����  � �          g� � �     b  ��  ��   ��  a       ���            �����  �  |         ����  � �          <x� � �     '  �  8B   ��  b       ��7            R  �  �  �         ����  � �          D~� � �     ^  ��  �W   ��  b       ��7            S  �  �  �         ����  � �          L�� � �     �  �  �l   ��  b       ��7            �����  �  �         ����  � �          k� �     �  ��  n
   ��  c       ��Y            (R  �  �  �         ����  � �          s��     &  V�  
7
   ��  c       ��Y            'S  �  �  �         ����  � �          {�
�     e  ��  �O
   ��  c       ��Y            &�����  �  �         ����  � �          ��2&�     X  ��  `>   ��  d       ��Z            5\  �  �  �         ����  � �          ��8,�     �  ��  �Z   ��  d       ��Z            4]  �  �  �         ����  � �          ��>2�     �  j�  �v   ��  d       ��Z            3�����  �  �         ����  e g          U� n b       )  X9        �       ��g            � 4  �  �  3         ����  q s          U� n b       )  X9        �       ��g            � 5  �  �  3         ����  � �          U� n b       )  X9        �       ��g            � �����  �  3         ����  m o          �� � �       �  �M  �   ��  �       ��h           	 � >  �  �  4         ����  z |          �� � �       �  O  <   ��  �       ��h           	 � ?  �  �  4         ����  � �          �� �         P  �    ��  �       ��h           	 � �����  �  4         ����  r t          �� �       J
  �]     ��  �     	  ��           
 � >  �  �           ����  � �          �$� �       k
  �^  �   ��  �     	  ��           
 � ?  �  �           ����  � �          �*� �       �
  �_  �   ��  �     	  ��           
 � �����  �           ����  z |          �=� � t     J  �n  �/   ��  �     
  ���            H  �  �  �         ����  � �          C� � u     r  �o  p?   ��  �     
  ���            I  �  �  �         ����  � �          I� � v     �  >q  �N   ��  �     
  ���            �����  �  �         ����   �          4[� � ~     �  L�  ܐ   ��  �       ���            H  �  �  ~         ����  � �          <a� �      �  ��  $�   ��  �       ���            I  �  �  ~         ����  � �          Dg� � �     .  �  l�   ��  �       ���            �����  �  ~         ����  � �          cx� � �     �  t�  X,   ��  �       ��<            R  �  �  �         ����  � �          k~� � �     &  ��  �A   ��  �       ��<            S  �  �  �         ����  � �          s�� � �     ]  ��   W   ��  �       ��<            �����  �  �         ����  � �          �� �     �  "�  �
   ��  �       ��e            (R  �  �  �         ����  � �          ���     �  Ƭ  �
   ��  �       ��e            'S  �  �  �         ����  � �          ��
�     )  j�  68
   ��  �       ��e            &�����  �  �         ����  � �          ��2&�       V�  `%   ��  �       ��f            5\  �  �  �         ����  � �          ��8,�     `  �  �A   ��  �       ��f            4]  �  �  �         ����  � �          ��>2�     �  ��  �]   ��  �       ��f            3�����  �  �         ����  c e          ;� n b         �7  �      )       ��z            � 4  �  �  F         ����  n q          ;� n b         �7  �      )       ��z            � 5  �  �  F         ����  ~ �          ;� n b         �7  �      )       ��z            � �����  �  F         ����  h j          �� � �       �  hL  �   ��  *     	  ��{           	 � >  �  �  G         ����  u w          �� � �       �  vM  �   ��  *     	  ��{           	 � ?  �  �  G         ����  � �          �� �       �  �N  (   ��  *     	  ��{           	 � �����  �  G         ����  p r          �� �       
  �[  ��   ��  +     
  ��           
 � >  �  �  
         ����  } �          �$� �       ?
  *]  �    ��  +     
  ��           
 � ?  �  �  
         ����  � �          �*� �       `
  V^  �   ��  +     
  ��           
 � �����  �  
         ����  v x          �=� � t       m  8   ��  ,       ���            H  �  �  �         ����  � �          �C� � u     B  dn  �,   ��  ,       ���            I  �  �  �         ����  � �          �I� � v     j  �o  (<   ��  ,       ���            �����  �  �         ����  ~           [� � ~     �  �  �|   ��  -       ���            H  �  �  }         ����  � �          "a� �      �  $�  Ԏ   ��  -       ���            I  �  �  }         ����  � �          *g� � �     �  ��  �   ��  -       ���            �����  �  }         ����  � �          Ix� � �     �  �  x   ��  .       ��A            R  �  �  �         ����  � �          Q~� � �     �  j�  �+   ��  .       ��A            S  �  �  �         ����  � �          Y�� � �     %  �   A   ��  .       ��A            �����  �  �         ����  � �          x� �     o  ��  ��	   ��  /       ��q            (R  �  �           ����  � �          ���     �  6�  *
   ��  /       ��q            'S  �  �           ����  � �          ��
�     �  ڬ  � 
   ��  /       ��q            &�����  �           ����  � �          ��2&�     �  ��  `   ��  0       ��r            5\  �  �           ����  � �          ��8,�        ��  �(   ��  0       ��r            4]  �  �           ����  � �          ��>2�     h  J�  �D   ��  0       ��r            3�����  �           ����  c e          M� n b       q  x<  8       �     �   �            � 4  �  �  Y         ����  n q          M� n b       q  x<  8       �     �   �            � 5  �  �  Y         ����  ~ �          M� n b       q  x<  8       �     �   �            � �����  �  Y         ����  j m          �� � �         Q  �*   ��  �     �   �           	 � >  �  �  Z         ����  w z          �� � �       7  &R  |5   ��  �     �   �           	 � ?  �  �  Z         ����  � �          �� �       R  4S  @   ��  �     �   �           	 � �����  �  Z         ����  p r          �� �       �
  �`  z'   ��  �     �   �           
 � >  �  �  �         ����  } �          �$� �       �
  �a  ^4   ��  �     �   �           
 � ?  �  �  �         ����  � �          �*� �       �
  c  BA   ��  �     �   �           
 � �����  �  �         ����  x z          �=� � t     �  �q  xU   ��  �     �   �            H  �  �  �         ����  � �          �C� � u     �  s  �d   ��  �     �   �            I  �  �  �         ����  � �          I� � v     �  ^t  ht   ��  �     �   �            �����  �  �         ����  ~           ,[� � ~     8  l�  |�   ��  �     �   �            H  �  �           ����  � �          4a� �      g  ԅ  ��   ��  �     �   �            I  �  �           ����  � �          <g� � �     �  <�  �   ��  �     �   �            �����  �           ����  � �          [x� � �     _  ��  X   ��  �     �   F            R  �  �  �         ����  � �          c~� � �     �  �  lm   ��  �     �   F            S  �  �  �         ����  � �          k�� � �     �  ��  ��   ��  �     �   F            �����  �  �         ����  � �          �� �     #  B�  �5
   ��  �     �   }            (R  �  �           ����  � �          ���     b  �  zN
   ��  �     �   }            'S  �  �           ����  � �          ��
�     �  ��  g
   ��  �     �   }            &�����  �           ����  � �          ��2&�     �  v�  `W   ��  �     �   ~            5\  �  �           ����  � �          ��8,�     �  8�  �s   ��  �     �   ~            4]  �  �           ����  � �          ��>2�     (   ��  ��   ��  �     �   ~            3�����  �           ����   U W          � � r�       {  �<  #   ��  1       ��            � 4  �  �  �          ����   ` a          � � y�       �  �=  x+   ��  1       ��            � 5  �  �  �          ����   m n          � � ��       �  �>  �3   ��  1       ��            � �����  �  �          ����   [ ]          � � ��       |  �J  p�   ��  2     	  ��           	 � >  �  �  �          ����   f h          �  ��       �  �K  ��   ��  2     	  ��           	 � ?  �  �  �          ����   t w          � ��       �  �L  �   ��  2     	  ��           	 � �����  �  �          ����   ` c          � ��       �	  nZ  ��   ��  3     
  ��           
 � >  �  �  �         ����   l n          � ��       
  �[  ��   ��  3     
  ��           
 � ?  �  �  �         ����   { ~          � ��       4
  �\  ��   ��  3     
  ��           
 � �����  �  �         ����   g h          � 8�� t     �  �k  x
   ��  4       ���            H  �  �  �         ����   s u          � >�� u       �l  �   ��  4       ���            I  �  �  �         ����   � �          � D�� v     :  n  h)   ��  4       ���            �����  �  �         ����   m o          W � ~     h  ,~  <h   ��  5       ���            H  �  �  �         ����   z |          ](�      �  �  �z   ��  5       ���            I  �  �  �         ����   � �          c0� �     �  ��  ̌   ��  5       ���            �����  �  �         ����   p r          uO� �       T�  �    ��  6       ��(            R  �  �  �         ����   } �          "{W� �     �  ړ  �   ��  6       ��(            S  �  �  �         ����   � �          '�_� �     �  `�  @+   ��  6       ��(            �����  �  �         ����   x z          D�~�     3  �  �	   ��  7       ��7            (R  �  �  �         ����   � �          J���     r  ��  ��	   ��  7       ��7            'S  �  �  �         ����   � �          P���     �  J�  V	
   ��  7       ��7            &�����  �  �         ����   ~           d��,�     �  6�  `�   ��  8       ��8            5\  �  �  �         ����   � �          j��2�     �  ��  �   ��  8       ��8            4]  �  �  �         ����   � �          p��8�     (  ��  �+   ��  8       ��8            3�����  �  �         ����  U W          � � ]�       N  �:  t   ��  �       ��             � 4  �  �  �          ����  ` a          � � d�       d  �;  �   ��  �       ��             � 5  �  �  �          ����  m n          � � k�       z  �<  T"   ��  �       ��             � �����  �  �          ����  [ ]          � � ��       J  �H  ��   ��  �     	  ��!           	 � >  �  �  �          ����  f h          � � ��       e  �I  t�   ��  �     	  ��!           	 � ?  �  �  �          ����  t w          � � ��       �   K   �   ��  �     	  ��!           	 � �����  �  �          ����  _ `          � � ��       �	  zX  >�   ��  �     
  ��	           
 � >  �  �  �         ����  k l          � ��       �	  �Y  "�   ��  �     
  ��	           
 � ?  �  �  �         ����  z {          � ��       �	  �Z  �   ��  �     
  ��	           
 � �����  �  �         ����  e g          � #�� t     �  �i  �   ��  �       ���            H  �  �  �         ����  q s          � )�� u     �  �j  �   ��  �       ���            I  �  �  �         ����  � �          � /�� v     �  *l  �   ��  �       ���            �����  �  �         ����  j m          � B� ~     '  8|  �N   ��  �       ���            H  �  �  �         ����  w z          � H�      V  �}   a   ��  �       ���            I  �  �  �         ����  � �          � N� �     �    hs   ��  �       ���            �����  �  �         ����  p r          `:� �     9  `�  @�   ��  �       ��-            R  �  �  �         ����  } �          fB� �     p  �  ��   ��  �       ��-            S  �  �  �         ����  � �          lJ� �     �  l�  �   ��  �       ��-            �����  �  �         ����  x z          /~i�     �  �  Һ	   ��  �       ��C            (R  �  �  �         ����  � �          5�q�     '  ��  n�	   ��  �       ��C            'S  �  �  �         ����  � �          ;�y�     f  V�  
�	   ��  �       ��C            &�����  �  �         ����  | ~          O��,�     H  B�   �   ��  �       ��D            5\  �  �  �         ����  � �          U��2�     �  �  @�   ��  �       ��D            4]  �  �  �         ����  � �          [��8�     �  ��  `   ��  �       ��D            3�����  �  �         ����  U W          � � j�       E  p:  �   ��         ��F            � 4  �  �           ����  ` a          � � q�       [  `;  `   ��         ��F            � 5  �  �           ����  m n          � � x�       q  P<  �   ��         ��F            � �����  �           ����  [ ]          � � ��       @  �H   �   ��  	     	  ��G           	 � >  �  �           ����  f h          � � ��       [  �I  ��   ��  	     	  ��G           	 � ?  �  �           ����  t w          � � ��       v  �J  �   ��  	     	  ��G           	 � �����  �           ����  _ `          � 
��       �	  X  ��   ��  
     
  ��           
 � >  �  �  �         ����  k l          � ��       �	  BY  ��   ��  
     
  ��           
 � ?  �  �  �         ����  z {          � ��       �	  nZ  ��   ��  
     
  ��           
 � �����  �  �         ����  e g          � 0�� t     �  2i  X�   ��         ���            H  �  �  �         ����  q s          � 6�� u     �  |j  ��   ��         ���            I  �  �  �         ����  � �          � <�� v     �  �k  H   ��         ���            �����  �  �         ����  j m          � O� ~       �{  �I   ��         ���            H  �  �  �         ����  w z          U �      I  <}  \   ��         ���            I  �  �  �         ����  � �          [(� �     x  �~  Tn   ��         ���            �����  �  �         ����  p r          mG� �     +  ��  ��   ��         ��3            R  �  �  �         ����  } �          sO� �     b  ��  �   ��         ��3            S  �  �  �         ����  � �          yW� �     �  �  p
   ��         ��3            �����  �  �         ����  x z          <�v�     �  ��  ��	   ��         ��O            (R  �  �  �         ����  � �          B�~�       N�  ��	   ��         ��O            'S  �  �  �         ����  � �          H���     W  �  .�	   ��         ��O            &�����  �  �         ����  | ~          \��,�     8  ޼  ��   ��         ��P            5\  �  �  �         ����  � �          b��2�     �  ��   �   ��         ��P            4]  �  �  �         ����  � �          h��8�     �  b�      ��         ��P            3�����  �  �         ����  U W          � � X�       �  xA  8M   ��  n       ��Y            � 4  �  �  %         ����  ` a          � � _�       �  hB  �U   ��  n       ��Y            � 5  �  �  %         ����  m n          � � f�         XC  ^   ��  n       ��Y            � �����  �  %         ����  [ ]          � � ��       �  �O  P   ��  o     	  ��Z           	 � >  �  �  &         ����  f h          � � ��         �P  �%   ��  o     	  ��Z           	 � ?  �  �  &         ����  t w          � � ��       *  �Q  h0   ��  o     	  ��Z           	 � �����  �  &         ����  _ `          � � ��       v
  _  J   ��  p     
  ��           
 � >  �  �            ����  k l          � � ��       �
  J`  .#   ��  p     
  ��           
 � ?  �  �            ����  z {          � ��       �
  va  0   ��  p     
  ��           
 � �����  �            ����  e g          � �� t     z  :p  �B   ��  q       ���            H  �  �  �         ����  q s          � $�� u     �  �q  0R   ��  q       ���            I  �  �  �         ����  � �          � *�� v     �  �r  �a   ��  q       ���            �����  �  �         ����  j m          � =� ~       ܂  ,�   ��  r       ���            H  �  �  �         ����  w z          � C�      3  D�  t�   ��  r       ���            I  �  �  �         ����  � �          � I� �     b  ��  ��   ��  r       ���            �����  �  �         ����  p r          [5� �     '  �  8B   ��  s       ��8            R  �  �  �         ����  } �          a=� �     ^  ��  �W   ��  s       ��8            S  �  �  �         ����  � �          gE� �     �  �  �l   ��  s       ��8            �����  �  �         ����  x z          *yd�     �  ��  n
   ��  t       ��[            (R  �  �  �         ����  � �          0l�     &  V�  
7
   ��  t       ��[            'S  �  �  �         ����  � �          6�t�     e  ��  �O
   ��  t       ��[            &�����  �  �         ����  | ~          J��,�     X  ��  `>   ��  u       ��\            5\  �  �  �         ����  � �          P��2�     �  ��  �Z   ��  u       ��\            4]  �  �  �         ����  � �          V��8�     �  j�  �v   ��  u       ��\            3�����  �  �         ����  U W          � � �       �  �?  (?   ��  �       ��l            � 4  �  �  8         ����  ` a          � � ��       �  �@  �G   ��  �       ��l            � 5  �  �  8         ����  m n          � � ��       �  �A  P   ��  �       ��l            � �����  �  8         ����  [ ]          � ��       �  �M  �   ��  �       ��m           	 � >  �  �  9         ����  f h          � ��       �  O  <   ��  �       ��m           	 � ?  �  �  9         ����  t w          � ��         P  �    ��  �       ��m           	 � �����  �  9         ����  ` c          � ��       J
  �]     ��  �     	  ��           
 � >  �  �           ����  l n          � $��       k
  �^  �   ��  �     	  ��           
 � ?  �  �           ����  { ~          � )��       �
  �_  �   ��  �     	  ��           
 � �����  �           ����  g h          � E�� t     J  �n  �/   ��  �     
  ���            H  �  �  �         ����  s u          � K�� u     r  �o  p?   ��  �     
  ���            I  �  �  �         ����  � �          Q� v     �  >q  �N   ��  �     
  ���            �����  �  �         ����  m o          d-� ~     �  L�  ܐ   ��  �       ���            H  �  �  �         ����  z |          j5�      �  ��  $�   ��  �       ���            I  �  �  �         ����  � �          p=� �     .  �  l�   ��  �       ���            �����  �  �         ����  p r          )�\� �     �  t�  X,   ��  �       ��=            R  �  �  �         ����  } �          .�d� �     &  ��  �A   ��  �       ��=            S  �  �  �         ����  � �          3�l� �     ]  ��   W   ��  �       ��=            �����  �  �         ����  x z          P���     �  "�  �
   ��  �       ��g            (R  �  �  �         ����  � �          V���     �  Ƭ  �
   ��  �       ��g            'S  �  �  �         ����  � �          \���     )  j�  68
   ��  �       ��g            &�����  �  �         ����  ~           p��,�       V�  `%   ��  �       ��h            5\  �  �  �         ����  � �          v��2�     `  �  �A   ��  �       ��h            4]  �  �  �         ����  � �          |��8�     �  ��  �]   ��  �       ��h            3�����  �  �         ����  U W          � � e�       �  X>  1   ��  :       ��            � 4  �  �  K         ����  ` a          � � l�       �  H?  �9   ��  :       ��            � 5  �  �  K         ����  m n          � � s�       �  8@  �A   ��  :       ��            � �����  �  K         ����  [ ]          � � ��       �  hL  �   ��  ;     	  ���           	 � >  �  �  L         ����  f h          � � ��       �  vM  �   ��  ;     	  ���           	 � ?  �  �  L         ����  t w          � � ��       �  �N  (   ��  ;     	  ���           	 � �����  �  L         ����  _ `          � ��       
  �[  ��   ��  <     
  ��!           
 � >  �  �           ����  k l          � 
��       ?
  *]  �    ��  <     
  ��!           
 � ?  �  �           ����  z {          � ��       `
  V^  �   ��  <     
  ��!           
 � �����  �           ����  e g          � +�� t       m  8   ��  =       ���            H  �  �  �         ����  q s          � 1�� u     B  dn  �,   ��  =       ���            I  �  �  �         ����  � �          � 7�� v     j  �o  (<   ��  =       ���            �����  �  �         ����  j m          � J� ~     �  �  �|   ��  >       ���            H  �  �  �         ����  w z          � P�      �  $�  Ԏ   ��  >       ���            I  �  �  �         ����  � �          V#� �     �  ��  �   ��  >       ���            �����  �  �         ����  p r          hB� �     �  �  x   ��  ?       ��B            R  �  �  �         ����  } �          nJ� �     �  j�  �+   ��  ?       ��B            S  �  �  �         ����  � �          tR� �     %  �   A   ��  ?       ��B            �����  �  �         ����  x z          7�q�     o  ��  ��	   ��  @       ��s            (R  �  �           ����  � �          =�y�     �  6�  *
   ��  @       ��s            'S  �  �           ����  � �          C���     �  ڬ  � 
   ��  @       ��s            &�����  �           ����  | ~          W��,�     �  ��  `   ��  A       ��t            5\  �  �           ����  � �          ]��2�        ��  �(   ��  A       ��t            4]  �  �           ����  � �          c��8�     h  J�  �D   ��  A       ��t            3�����  �           ����  U W          � � w�         C  H[   ��  �     �   �            � 4  �  �  ^         ����  ` a          � � ~�       !  �C  �c   ��  �     �   �            � 5  �  �  ^         ����  m n          � � ��       7  �D  (l   ��  �     �   �            � �����  �  ^         ����  [ ]          �  ��         Q  �*   ��  �     �   �           	 � >  �  �  _         ����  f h          � ��       7  &R  |5   ��  �     �   �           	 � ?  �  �  _         ����  t w          � 
��       R  4S  @   ��  �     �   �           	 � �����  �  _         ����  ` c          � ��       �
  �`  z'   ��  �     �   �           
 � >  �  �  �         ����  l n          � ��       �
  �a  ^4   ��  �     �   �           
 � ?  �  �  �         ����  { ~          � !��       �
  c  BA   ��  �     �   �           
 � �����  �  �         ����  g h          � =�� t     �  �q  xU   ��  �     �   �            H  �  �  �         ����  s u          � C�� u     �  s  �d   ��  �     �   �            I  �  �  �         ����  � �          � I�� v     �  ^t  ht   ��  �     �   �            �����  �  �         ����  m o          
\%� ~     8  l�  |�   ��  �     �   �            H  �  �  �         ����  z |          b-�      g  ԅ  ��   ��  �     �   �            I  �  �  �         ����  � �          h5� �     �  <�  �   ��  �     �   �            �����  �  �         ����  p r          !zT� �     _  ��  X   ��  �     �   G            R  �  �  �         ����  } �          &�\� �     �  �  lm   ��  �     �   G            S  �  �  �         ����  � �          +�d� �     �  ��  ��   ��  �     �   G            �����  �  �         ����  x z          H���     #  B�  �5
   ��  �     �               (R  �  �           ����  � �          N���     b  �  zN
   ��  �     �               'S  �  �           ����  � �          T���     �  ��  g
   ��  �     �               &�����  �           ����  ~           h��,�     �  v�  `W   ��  �     �   �            5\  �  �           ����  � �          n��2�     �  8�  �s   ��  �     �   �            4]  �  �           ����  � �          t��8�     (   ��  ��   ��  �     �   �            3�����  �           ����   U W          6} 6       {  �<  #   ��  E       ��            � 4  �  �  �          ����   ` a          <� <�       �  �=  x+   ��  E       ��            � 5  �  �  �          ����   m n          B� B�       �  �>  �3   ��  E       ��            � �����  �  �          ����   [ ]          V� V�       |  �J  p�   ��  F     	  ��           	 � >  �  �  �          ����   f h          \� \�       �  �K  ��   ��  F     	  ��           	 � ?  �  �  �          ����   t w          b� b�       �  �L  �   ��  F     	  ��           	 � �����  �  �          ����   _ `          v� v�       �	  nZ  ��   ��  G     
  ��           
 � >  �  �  �         ����   k l          |� |�       
  �[  ��   ��  G     
  ��           
 � ?  �  �  �         ����   z {          �� ��       4
  �\  ��   ��  G     
  ��           
 � �����  �  �         ����   e g          �� �� t     �  �k  x
   ��  H       ���            H  �  �  �         ����   q s          �� �� u       �l  �   ��  H       ���            I  �  �  �         ����   � �          �� �� v     :  n  h)   ��  H       ���            �����  �  �         ����   j m          �� �� ~     h  ,~  <h   ��  I       ���            H  �  �  �         ����   w z          �� ��      �  �  �z   ��  I       ���            I  �  �  �         ����   � �          �� �� �     �  ��  ̌   ��  I       ���            �����  �  �         ����   p r          �� �� �       T�  �    ��  J       ��)            R  �  �  �         ����   } �          �� �� �     �  ړ  �   ��  J       ��)            S  �  �  �         ����   � �          � � �     �  `�  @+   ��  J       ��)            �����  �  �         ����   x z          � �     3  �  �	   ��  K       ��9            (R  �  �  �         ����   � �          ""�     r  ��  ��	   ��  K       ��9            'S  �  �  �         ����   � �          )	)�     �  J�  V	
   ��  K       ��9            &�����  �  �         ����   | ~          Q%Q'�     �  6�  `�   ��  L       ��:            5\  �  �  �         ����   � �          Y+Y-�     �  ��  �   ��  L       ��:            4]  �  �  �         ����   � �          a1a3�     (  ��  �+   ��  L       ��:            3�����  �  �         ����  S U          !} !       N  �:  t   ��  �       ��)            � 4  �  �  �          ����  ] `          '� '�       d  �;  �   ��  �       ��)            � 5  �  �  �          ����  j m          -� -�       z  �<  T"   ��  �       ��)            � �����  �  �          ����  Y [          A� A�       J  �H  ��   ��  �     	  ��*           	 � >  �  �  �          ����  c f          G� G�       e  �I  t�   ��  �     	  ��*           	 � ?  �  �  �          ����  q t          M� M�       �   K   �   ��  �     	  ��*           	 � �����  �  �          ����  _ `          a� a�       �	  zX  >�   ��  �     
  ��           
 � >  �  �  �         ����  k l          g� g�       �	  �Y  "�   ��  �     
  ��           
 � ?  �  �  �         ����  z {          m� m�       �	  �Z  �   ��  �     
  ��           
 � �����  �  �         ����  c e          �� �� t     �  �i  �   ��  �       ���            H  �  �  �         ����  n q          �� �� u     �  �j  �   ��  �       ���            I  �  �  �         ����  ~ �          �� �� v     �  *l  �   ��  �       ���            �����  �  �         ����  h j          �� �� ~     '  8|  �N   ��  �       ���            H  �  �  �         ����  u w          �� ��      V  �}   a   ��  �       ���            I  �  �  �         ����  � �          �� �� �     �    hs   ��  �       ���            �����  �  �         ����  o p          �� �� �     9  `�  @�   ��  �       ��.            R  �  �  �         ����  | }          �� �� �     p  �  ��   ��  �       ��.            S  �  �  �         ����  � �          �� �� �     �  l�  �   ��  �       ��.            �����  �  �         ����  v x          � �     �  �  Һ	   ��  �       ��E            (R  �  �  �         ����  � �          �     '  ��  n�	   ��  �       ��E            'S  �  �  �         ����  � �          	�     f  V�  
�	   ��  �       ��E            &�����  �  �         ����  | ~          <%<'�     H  B�   �   ��  �       ��F            5\  �  �  �         ����  � �          D+D-�     �  �  @�   ��  �       ��F            4]  �  �  �         ����  � �          L1L3�     �  ��  `   ��  �       ��F            3�����  �  �         ����  S U          .} .       E  p:  �   ��         ��O            � 4  �  �           ����  ] `          4� 4�       [  `;  `   ��         ��O            � 5  �  �           ����  j m          :� :�       q  P<  �   ��         ��O            � �����  �           ����  Y [          N� N�       @  �H   �   ��       	  ��P           	 � >  �  �           ����  c f          T� T�       [  �I  ��   ��       	  ��P           	 � ?  �  �           ����  q t          Z� Z�       v  �J  �   ��       	  ��P           	 � �����  �           ����  _ `          n� n�       �	  X  ��   ��       
  ��           
 � >  �  �  �         ����  k l          t� t�       �	  BY  ��   ��       
  ��           
 � ?  �  �  �         ����  z {          z� z�       �	  nZ  ��   ��       
  ��           
 � �����  �  �         ����  c e          �� �� t     �  2i  X�   ��         ���            H  �  �  �         ����  n q          �� �� u     �  |j  ��   ��         ���            I  �  �  �         ����  ~ �          �� �� v     �  �k  H   ��         ���            �����  �  �         ����  h j          �� �� ~       �{  �I   ��         ���            H  �  �  �         ����  u w          �� ��      I  <}  \   ��         ���            I  �  �  �         ����  � �          �� �� �     x  �~  Tn   ��         ���            �����  �  �         ����  o p          �� �� �     +  ��  ��   ��         ��4            R  �  �  �         ����  | }          �� �� �     b  ��  �   ��         ��4            S  �  �  �         ����  � �          �� �� �     �  �  p
   ��         ��4            �����  �  �         ����  v x          � �     �  ��  ��	   ��         ��Q            (R  �  �  �         ����  � �          �       N�  ��	   ��         ��Q            'S  �  �  �         ����  � �          !	!�     W  �  .�	   ��         ��Q            &�����  �  �         ����  | ~          I%I'�     8  ޼  ��   ��          ��R            5\  �  �  �         ����  � �          Q+Q-�     �  ��   �   ��          ��R            4]  �  �  �         ����  � �          Y1Y3�     �  b�      ��          ��R            3�����  �  �         ����  S U          }        �  xA  8M   ��         ��b            � 4  �  �  .         ����  ] `          "� "�       �  hB  �U   ��         ��b            � 5  �  �  .         ����  j m          (� (�         XC  ^   ��         ��b            � �����  �  .         ����  Y [          <� <�       �  �O  P   ��  �     	  ��c           	 � >  �  �  /         ����  c f          B� B�         �P  �%   ��  �     	  ��c           	 � ?  �  �  /         ����  q t          H� H�       *  �Q  h0   ��  �     	  ��c           	 � �����  �  /         ����  _ `          \� \�       v
  _  J   ��  �     
  ��           
 � >  �  �           ����  k l          b� b�       �
  J`  .#   ��  �     
  ��           
 � ?  �  �           ����  z {          h� h�       �
  va  0   ��  �     
  ��           
 � �����  �           ����  c e          �� �� t     z  :p  �B   ��  �       ���            H  �  �  �         ����  n q          �� �� u     �  �q  0R   ��  �       ���            I  �  �  �         ����  ~ �          �� �� v     �  �r  �a   ��  �       ���            �����  �  �         ����  h j          �� �� ~       ܂  ,�   ��  �       ���            H  �  �  �         ����  u w          �� ��      3  D�  t�   ��  �       ���            I  �  �  �         ����  � �          �� �� �     b  ��  ��   ��  �       ���            �����  �  �         ����  o p          �� �� �     '  �  8B   ��  �       ��9            R  �  �  �         ����  | }          �� �� �     ^  ��  �W   ��  �       ��9            S  �  �  �         ����  � �          �� �� �     �  �  �l   ��  �       ��9            �����  �  �         ����  v x          � �     �  ��  n
   ��  �       ��]            (R  �  �  �         ����  � �          �     &  V�  
7
   ��  �       ��]            'S  �  �  �         ����  � �          	�     e  ��  �O
   ��  �       ��]            &�����  �  �         ����  | ~          7%7'�     X  ��  `>   ��  �       ��^            5\  �  �  �         ����  � �          ?+?-�     �  ��  �Z   ��  �       ��^            4]  �  �  �         ����  � �          G1G3�     �  j�  �v   ��  �       ��^            3�����  �  �         ����  U W          C} C       �  �?  (?   ��  �       ��u            � 4  �  �  A         ����  ` a          I� I�       �  �@  �G   ��  �       ��u            � 5  �  �  A         ����  m n          O� O�       �  �A  P   ��  �       ��u            � �����  �  A         ����  [ ]          c� c�       �  �M  �   ��  �       ��v           	 � >  �  �  B         ����  f h          i� i�       �  O  <   ��  �       ��v           	 � ?  �  �  B         ����  t w          o� o�         P  �    ��  �       ��v           	 � �����  �  B         ����  _ `          �� ��       J
  �]     ��  �     	  ��           
 � >  �  �           ����  k l          �� ��       k
  �^  �   ��  �     	  ��           
 � ?  �  �           ����  z {          �� ��       �
  �_  �   ��  �     	  ��           
 � �����  �           ����  e g          �� �� t     J  �n  �/   ��  �     
  ���            H  �  �  �         ����  q s          �� �� u     r  �o  p?   ��  �     
  ���            I  �  �  �         ����  � �          �� �� v     �  >q  �N   ��  �     
  ���            �����  �  �         ����  j m          �� �� ~     �  L�  ܐ   ��  �       ���            H  �  �  �         ����  w z          �� ��      �  ��  $�   ��  �       ���            I  �  �  �         ����  � �          �� �� �     .  �  l�   ��  �       ���            �����  �  �         ����  p r          � � �     �  t�  X,   ��  �       ��>            R  �  �  �         ����  } �          � � �     &  ��  �A   ��  �       ��>            S  �  �  �         ����  � �          � � �     ]  ��   W   ��  �       ��>            �����  �  �         ����  x z          (� (�     �  "�  �
   ��  �       ��i            (R  �  �  �         ����  � �          //�     �  Ƭ  �
   ��  �       ��i            'S  �  �  �         ����  � �          6	6�     )  j�  68
   ��  �       ��i            &�����  �  �         ����  | ~          ^%^'�       V�  `%   ��  �       ��j            5\  �  �  �         ����  � �          f+f-�     `  �  �A   ��  �       ��j            4]  �  �  �         ����  � �          n1n3�     �  ��  �]   ��  �       ��j            3�����  �  �         ����  S U          )} )       �  X>  1   ��  K       ���            � 4  �  �  T         ����  ] `          /� /�       �  H?  �9   ��  K       ���            � 5  �  �  T         ����  j m          5� 5�       �  8@  �A   ��  K       ���            � �����  �  T         ����  Y [          I� I�       �  hL  �   ��  L     	  ���           	 � >  �  �  U         ����  c f          O� O�       �  vM  �   ��  L     	  ���           	 � ?  �  �  U         ����  q t          U� U�       �  �N  (   ��  L     	  ���           	 � �����  �  U         ����  _ `          i� i�       
  �[  ��   ��  M     
  ��#           
 � >  �  �           ����  k l          o� o�       ?
  *]  �    ��  M     
  ��#           
 � ?  �  �           ����  z {          u� u�       `
  V^  �   ��  M     
  ��#           
 � �����  �           ����  c e          �� �� t       m  8   ��  N       ���            H  �  �  �         ����  n q          �� �� u     B  dn  �,   ��  N       ���            I  �  �  �         ����  ~ �          �� �� v     j  �o  (<   ��  N       ���            �����  �  �         ����  h j          �� �� ~     �  �  �|   ��  O       ���            H  �  �  �         ����  u w          �� ��      �  $�  Ԏ   ��  O       ���            I  �  �  �         ����  � �          �� �� �     �  ��  �   ��  O       ���            �����  �  �         ����  o p          �� �� �     �  �  x   ��  P       ��C            R  �  �  �         ����  | }          �� �� �     �  j�  �+   ��  P       ��C            S  �  �  �         ����  � �          �� �� �     %  �   A   ��  P       ��C            �����  �  �         ����  v x          � �     o  ��  ��	   ��  Q       ��u            (R  �  �           ����  � �          �     �  6�  *
   ��  Q       ��u            'S  �  �           ����  � �          	�     �  ڬ  � 
   ��  Q       ��u            &�����  �           ����  x z          D%D'�     �  ��  `   ��  R       ��v            5\  �  �  	         ����  � �          L+L-�        ��  �(   ��  R       ��v            4]  �  �  	         ����  � �          T1T3�     h  J�  �D   ��  R       ��v            3�����  �  	         ����  U W          ;} ;         C  H[   ��  �     �   �            � 4  �  �  g         ����  ` a          A� A�       !  �C  �c   ��  �     �   �            � 5  �  �  g         ����  m n          G� G�       7  �D  (l   ��  �     �   �            � �����  �  g         ����  [ ]          [� [�         Q  �*   ��  �     �   �           	 � >  �  �  h         ����  f h          a� a�       7  &R  |5   ��  �     �   �           	 � ?  �  �  h         ����  t w          g� g�       R  4S  @   ��  �     �   �           	 � �����  �  h         ����  _ `          {� {�       �
  �`  z'   ��  �     �   �           
 � >  �  �  �         ����  k l          �� ��       �
  �a  ^4   ��  �     �   �           
 � ?  �  �  �         ����  z {          �� ��       �
  c  BA   ��  �     �   �           
 � �����  �  �         ����  e g          �� �� t     �  �q  xU   ��  �     �   �            H  �  �  �         ����  q s          �� �� u     �  s  �d   ��  �     �   �            I  �  �  �         ����  � �          �� �� v     �  ^t  ht   ��  �     �   �            �����  �  �         ����  j m          �� �� ~     8  l�  |�   ��  �     �   �            H  �  �  �         ����  w z          �� ��      g  ԅ  ��   ��  �     �   �            I  �  �  �         ����  � �          �� �� �     �  <�  �   ��  �     �   �            �����  �  �         ����  p r          �� �� �     _  ��  X   ��  �     �   H            R  �  �  �         ����  } �           �  � �     �  �  lm   ��  �     �   H            S  �  �  �         ����  � �          � � �     �  ��  ��   ��  �     �   H            �����  �  �         ����  x z           �  �     #  B�  �5
   ��  �     �   �            (R  �  �           ����  � �          ''�     b  �  zN
   ��  �     �   �            'S  �  �           ����  � �          .	.�     �  ��  g
   ��  �     �   �            &�����  �           ����  | ~          V%V'�     �  v�  `W   ��  �     �   �            5\  �  �           ����  � �          ^+^-�     �  8�  �s   ��  �     �   �            4]  �  �           ����  � �          f1f3�     (   ��  ��   ��  �     �   �            3�����  �           ����   I L          � � t�       {  �<  #   ��  Y       ��(            � 4  �  �           ����   R U          � � {�       �  �=  x+   ��  Y       ��(            � 5  �  �           ����   ^ `          � � ��       �  �>  �3   ��  Y       ��(            � �����  �           ����   N O          � � ��       |  �J  p�   ��  Z     	  ��)           	 � >  �  �           ����   W X          � � ��       �  �K  ��   ��  Z     	  ��)           	 � ?  �  �           ����   c e          � � ��       �  �L  �   ��  Z     	  ��)           	 � �����  �           ����   Q S          � ��       �	  nZ  ��   ��  [     
  ��*           
 � >  �  �           ����   [ ]          � ��       
  �[  ��   ��  [     
  ��*           
 � ?  �  �           ����   g j          � ��       4
  �\  ��   ��  [     
  ��*           
 � �����  �           ����   W Y          � -�� t     �  �k  x
   ��  \       ���            H  �  �  �         ����   a c          � 3�� u       �l  �   ��  \       ���            I  �  �  �         ����   n q          � 9�� v     :  n  h)   ��  \       ���            �����  �  �         ����   [ ]          � L"� ~     h  ,~  <h   ��  ]       ���            H  �  �  �         ����   f h          � R*�      �  �  �z   ��  ]       ���            I  �  �  �         ����   t w          � X2� �     �  ��  ̌   ��  ]       ���            �����  �  �         ����   _ `          jQ� �       T�  �    ��  ^       ��*            R  �  �  �         ����   k l          pY� �     �  ړ  �   ��  ^       ��*            S  �  �  �         ����   z {          va� �     �  `�  @+   ��  ^       ��*            �����  �  �         ����   e g          /���     3  �  �	   ��  _       ��;            (R  �  �  �         ����   q s          5���     r  ��  ��	   ��  _       ��;            'S  �  �  �         ����   � �          ;���     �  J�  V	
   ��  _       ��;            &�����  �  �         ����   h j          O��-�     �  6�  `�   ��  `       ��<            5\  �  �  �         ����   u w          U��3�     �  ��  �   ��  `       ��<            4]  �  �  �         ����   � �          [��9�     (  ��  �+   ��  `       ��<            3�����  �  �         ����  I L          � � k|       N  �:  t   ��  �       ��-            � 4  �  �           ����  R U          � � r�       d  �;  �   ��  �       ��-            � 5  �  �           ����  ^ `          � � y�       z  �<  T"   ��  �       ��-            � �����  �           ����  N O          � � ��       J  �H  ��   ��  �     	  ��.           	 � >  �  �           ����  W X          � � ��       e  �I  t�   ��  �     	  ��.           	 � ?  �  �           ����  c e          � � ��       �   K   �   ��  �     	  ��.           	 � �����  �           ����  Q S          � � ��       �	  zX  >�   ��  �     
  ��/           
 � >  �  �           ����  [ ]          � ��       �	  �Y  "�   ��  �     
  ��/           
 � ?  �  �           ����  g j          � ��       �	  �Z  �   ��  �     
  ��/           
 � �����  �           ����  U W          � $�� t     �  �i  �   ��  �       ���            H  �  �  �         ����  ` a          � *�� u     �  �j  �   ��  �       ���            I  �  �  �         ����  m n          � 0�� v     �  *l  �   ��  �       ���            �����  �  �         ����  Y [          � C� ~     '  8|  �N   ��  �       ���            H  �  �  �         ����  c f          � I!�      V  �}   a   ��  �       ���            I  �  �  �         ����  q t          � O)� �     �    hs   ��  �       ���            �����  �  �         ����  ] _          � aH� �     9  `�  @�   ��  �       ��/            R  �  �  �         ����  h k          gP� �     p  �  ��   ��  �       ��/            S  �  �  �         ����  w z          	mX� �     �  l�  �   ��  �       ��/            �����  �  �         ����  c e          &w� �     �  �  Һ	   ��  �       ��G            (R  �  �  �         ����  n q          ,��     '  ��  n�	   ��  �       ��G            'S  �  �  �         ����  ~ �          2���     f  V�  
�	   ��  �       ��G            &�����  �  �         ����  g h          F��$�     H  B�   �   ��  �       ��H            5\  �  �  �         ����  s u          L��*�     �  �  @�   ��  �       ��H            4]  �  �  �         ����  � �          R��0�     �  ��  `   ��  �       ��H            3�����  �  �         ����  I L          � � n�       E  p:  �   ��  *       ��2            � 4  �  �           ����  R U          � � u�       [  `;  `   ��  *       ��2            � 5  �  �           ����  ^ `          � � |�       q  P<  �   ��  *       ��2            � �����  �           ����  N O          � � ��       @  �H   �   ��  +     	  ��3           	 � >  �  �           ����  W X          � � ��       [  �I  ��   ��  +     	  ��3           	 � ?  �  �           ����  c e          � � ��       v  �J  �   ��  +     	  ��3           	 � �����  �           ����  Q S          � 	��       �	  X  ��   ��  ,     
  ��4           
 � >  �  �           ����  [ ]          � ��       �	  BY  ��   ��  ,     
  ��4           
 � ?  �  �           ����  g j          � ��       �	  nZ  ��   ��  ,     
  ��4           
 � �����  �           ����  U W          � /�� t     �  2i  X�   ��  -       ���            H  �  �  �         ����  ` a          � 5�� u     �  |j  ��   ��  -       ���            I  �  �  �         ����  m n          � ;�� v     �  �k  H   ��  -       ���            �����  �  �         ����  Y [          � N� ~       �{  �I   ��  .       ���            H  �  �  �         ����  c f          � T$�      I  <}  \   ��  .       ���            I  �  �  �         ����  q t          Z,� �     x  �~  Tn   ��  .       ���            �����  �  �         ����  ] _          lK� �     +  ��  ��   ��  /       ��5            R  �  �  �         ����  h k          rS� �     b  ��  �   ��  /       ��5            S  �  �  �         ����  w z          x[� �     �  �  p
   ��  /       ��5            �����  �  �         ����  c e          8�z�     �  ��  ��	   ��  0       ��S            (R  �  �  �         ����  n q          >���       N�  ��	   ��  0       ��S            'S  �  �  �         ����  ~ �          D���     W  �  .�	   ��  0       ��S            &�����  �  �         ����  g h          X��-�     8  ޼  ��   ��  1       ��T            5\  �  �  �         ����  s u          ^��3�     �  ��   �   ��  1       ��T            4]  �  �  �         ����  � �          d��9�     �  b�      ��  1       ��T            3�����  �  �         ����  I L          � � hy       �  xA  8M   ��  �       ��7            � 4  �  �  !         ����  R U          � � o}       �  hB  �U   ��  �       ��7            � 5  �  �  !         ����  ^ `          � � v�         XC  ^   ��  �       ��7            � �����  �  !         ����  N O          � � ��       �  �O  P   ��  �     	  ��8           	 � >  �  �  "         ����  W X          � � ��         �P  �%   ��  �     	  ��8           	 � ?  �  �  "         ����  c e          � � ��       *  �Q  h0   ��  �     	  ��8           	 � �����  �  "         ����  Q S          � � ��       v
  _  J   ��  �     
  ��9           
 � >  �  �  #         ����  [ ]          �  ��       �
  J`  .#   ��  �     
  ��9           
 � ?  �  �  #         ����  g j          � ��       �
  va  0   ��  �     
  ��9           
 � �����  �  #         ����  U W          � !�� t     z  :p  �B   ��  �       ���            H  �  �  �         ����  ` a          � '�� u     �  �q  0R   ��  �       ���            I  �  �  �         ����  m n          � -�� v     �  �r  �a   ��  �       ���            �����  �  �         ����  Y [          � @� ~       ܂  ,�   ��  �       ���            H  �  �  �         ����  c f          � F�      3  D�  t�   ��  �       ���            I  �  �  �         ����  q t          � L&� �     b  ��  ��   ��  �       ���            �����  �  �         ����  ] _          � ^E� �     '  �  8B   ��  �       ��:            R  �  �  �         ����  h k          dM� �     ^  ��  �W   ��  �       ��:            S  �  �  �         ����  w z          jU� �     �  �  �l   ��  �       ��:            �����  �  �         ����  c e          #|t� �     �  ��  n
   ��  �       ��_            (R  �  �  �         ����  n q          )�| �     &  V�  
7
   ��  �       ��_            'S  �  �  �         ����  ~ �          /���     e  ��  �O
   ��  �       ��_            &�����  �  �         ����  g h          C��!�     X  ��  `>   ��  �       ��`            5\  �  �  �         ����  s u          I��'�     �  ��  �Z   ��  �       ��`            4]  �  �  �         ����  � �          O��-�     �  j�  �v   ��  �       ��`            3�����  �  �         ����  I L          � � ��       �  �?  (?   ��  �       ��<            � 4  �  �  &         ����  R U          � � ��       �  �@  �G   ��  �       ��<            � 5  �  �  &         ����  ^ `          � � ��       �  �A  P   ��  �       ��<            � �����  �  &         ����  N O          � � ��       �  �M  �   ��  �       ��=           	 � >  �  �  '         ����  W X          � ��       �  O  <   ��  �       ��=           	 � ?  �  �  '         ����  c e          � 	��         P  �    ��  �       ��=           	 � �����  �  '         ����  Q S          � ��       J
  �]     ��  �     	  ��>           
 � >  �  �  (         ����  [ ]          � ��       k
  �^  �   ��  �     	  ��>           
 � ?  �  �  (         ����  g j          �  ��       �
  �_  �   ��  �     	  ��>           
 � �����  �  (         ����  W Y          � <�� t     J  �n  �/   ��  �     
  ���            H  �  �  �         ����  a c          � B� u     r  �o  p?   ��  �     
  ���            I  �  �  �         ����  n q          � H	� v     �  >q  �N   ��  �     
  ���            �����  �  �         ����  [ ]           [1� ~     �  L�  ܐ   ��  �       ���            H  �  �  �         ����  f h          a9�      �  ��  $�   ��  �       ���            I  �  �  �         ����  t w          
gA� �     .  �  l�   ��  �       ���            �����  �  �         ����  _ `          y`� �     �  t�  X,   ��  �       ��?            R  �  �  �         ����  k l          h�     &  ��  �A   ��  �       ��?            S  �  �  �         ����  z {          !�p	�     ]  ��   W   ��  �       ��?            �����  �  �         ����  e g          >���     �  "�  �
   ��  �       ��k            (R  �  �  �         ����  q s          D���     �  Ƭ  �
   ��  �       ��k            'S  �  �  �         ����  � �          J�� �     )  j�  68
   ��  �       ��k            &�����  �  �         ����  h j          ^��<�       V�  `%   ��  �       ��l            5\  �  �  �         ����  u w          d��B�     `  �  �A   ��  �       ��l            4]  �  �  �         ����  � �          j��H�     �  ��  �]   ��  �       ��l            3�����  �  �         ����  I L          � � z�       �  X>  1   ��  \       ��A            � 4  �  �  +         ����  R U          � � ��       �  H?  �9   ��  \       ��A            � 5  �  �  +         ����  ^ `          � � ��       �  8@  �A   ��  \       ��A            � �����  �  +         ����  N O          � � ��       �  hL  �   ��  ]     	  ��B           	 � >  �  �  ,         ����  W X          � � ��       �  vM  �   ��  ]     	  ��B           	 � ?  �  �  ,         ����  c e          �  ��       �  �N  (   ��  ]     	  ��B           	 � �����  �  ,         ����  Q S          � ��       
  �[  ��   ��  ^     
  ��C           
 � >  �  �  -         ����  [ ]          � ��       ?
  *]  �    ��  ^     
  ��C           
 � ?  �  �  -         ����  g j          � ��       `
  V^  �   ��  ^     
  ��C           
 � �����  �  -         ����  U W          � 3�� t       m  8   ��  _       ���            H  �  �  �         ����  ` a          � 9�� u     B  dn  �,   ��  _       ���            I  �  �  �         ����  m n          � ? � v     j  �o  (<   ��  _       ���            �����  �  �         ����  Y [          � R(� ~     �  �  �|   ��  `       ���            H  �  �  �         ����  c f          � X0�      �  $�  Ԏ   ��  `       ���            I  �  �  �         ����  q t          ^8� �     �  ��  �   ��  `       ���            �����  �  �         ����  ] _          pW� �     �  �  x   ��  a       ��D            R  �  �  �         ����  h k          v_� �     �  j�  �+   ��  a       ��D            S  �  �  �         ����  w z          |g �     %  �   A   ��  a       ��D            �����  �  �         ����  c e          5���     o  ��  ��	   ��  b       ��w            (R  �  �  
         ����  n q          ;���     �  6�  *
   ��  b       ��w            'S  �  �  
         ����  ~ �          A���     �  ڬ  � 
   ��  b       ��w            &�����  �  
         ����  g h          U��3�     �  ��  `   ��  c       ��x            5\  �  �           ����  s u          [��9�        ��  �(   ��  c       ��x            4]  �  �           ����  � �          a��?�     h  J�  �D   ��  c       ��x            3�����  �           ����  L N          � � b�         C  H[   ��  �     �   �            � 4  �  �  �         ����  U W          � � i�       !  �C  �c   ��  �     �   �            � 5  �  �  �         ����  ` c          � � p�       7  �D  (l   ��  �     �   �            � �����  �  �         ����  O Q          � � ��         Q  �*   ��  �     �   �           	 � >  �  �  �         ����  X [          � � ��       7  &R  |5   ��  �     �   �           	 � ?  �  �  �         ����  e g          � � ��       R  4S  @   ��  �     �   �           	 � �����  �  �         ����  S U          � � ��       �
  �`  z'   ��  �     �   �           
 � >  �  �  �         ����  ] `          � � ��       �
  �a  ^4   ��  �     �   �           
 � ?  �  �  �         ����  j m          � ��       �
  c  BA   ��  �     �   �           
 � �����  �  �         ����  W Y          �  �� t     �  �q  xU   ��  �     �   �            H  �  �  �         ����  a c          � &�� u     �  s  �d   ��  �     �   �            I  �  �  �         ����  n q          � ,�� v     �  ^t  ht   ��  �     �   �            �����  �  �         ����  [ ]          � ?� ~     8  l�  |�   ��  �     �   �            H  �  �  �         ����  f h          � E�      g  ԅ  ��   ��  �     �   �            I  �  �  �         ����  t w          � K � �     �  <�  �   ��  �     �   �            �����  �  �         ����  _ `          ]?� �     _  ��  X   ��  �     �   I            R  �  �  �         ����  k l          
cG� �     �  �  lm   ��  �     �   I            S  �  �  �         ����  z {          iO� �     �  ��  ��   ��  �     �   I            �����  �  �         ����  g h          ,{n�     #  B�  �5
   ��  �     �   �            (R  �  �           ����  s u          2�v	�     b  �  zN
   ��  �     �   �            'S  �  �           ����  � �          8�~�     �  ��  g
   ��  �     �   �            &�����  �           ����  j m          L��*�     �  v�  `W   ��  �     �   �            5\  �  �           ����  w z          R��0�     �  8�  �s   ��  �     �   �            4]  �  �           ����  � �          X��6�     (   ��  ��   ��  �     �   �            3�����  �           ����   U W          )� ~       {  �<  #   ��  m       ��}            � 4  �  �  =         ����   ` a           /� �       �  �=  x+   ��  m       ��}            � 5  �  �  =         ����   m n          &5� �       �  �>  �3   ��  m       ��}            � �����  �  =         ����   [ ]          :H� �       |  �J  p�   ��  n     	  ���           	 � >  �  �  I         ����   f h          @N� �       �  �K  ��   ��  n     	  ���           	 � ?  �  �  I         ����   t w          FT� �       �  �L  �   ��  n     	  ���           	 � �����  �  I         ����   ` c          Zf� �       �	  nZ  ��   ��  o     
  ���           
 � >  �  �  U         ����   l n          `l� �       
  �[  ��   ��  o     
  ���           
 � ?  �  �  U         ����   { ~          fr� �       4
  �\  ��   ��  o     
  ���           
 � �����  �  U         ����   g h          ��� � t     �  �k  x
   ��  p       ���            H  �  �  a         ����   s u          ��� � u       �l  �   ��  p       ���            I  �  �  a         ����   � �          ��� � v     :  n  h)   ��  p       ���            �����  �  a         ����   m o          ��� � ~     h  ,~  <h   ��  q       ���            H  �  �  m         ����   z |          ��� �      �  �  �z   ��  q       ���            I  �  �  m         ����   � �          ��� � �     �  ��  ̌   ��  q       ���            �����  �  m         ����   p r          ��� � �       T�  �    ��  r       ��+            R  �  �  �         ����   } �          ��� � �     �  ړ  �   ��  r       ��+            S  �  �  �         ����   � �          ��� � �     �  `�  @+   ��  r       ��+            �����  �  �         ����   x z          � �     3  �  �	   ��  s       ��=            (R  �  �  �         ����   � �          
�     r  ��  ��	   ��  s       ��=            'S  �  �  �         ����   � �          
�     �  J�  V	
   ��  s       ��=            &�����  �  �         ����   ~           572&�     �  6�  `�   ��  t       ��>            5\  �  �  �         ����   � �          =?8,�     �  ��  �   ��  t       ��>            4]  �  �  �         ����   � �          EG>2�     (  ��  �+   ��  t       ��>            3�����  �  �         ����  U W          � ~       N  �:  t   ��  �       ��            � 4  �  �  ?         ����  ` a           %� �       d  �;  �   ��  �       ��            � 5  �  �  ?         ����  m n          &+� �       z  �<  T"   ��  �       ��            � �����  �  ?         ����  [ ]          :>� �       J  �H  ��   ��  �     	  ���           	 � >  �  �  K         ����  f h          @D� �       e  �I  t�   ��  �     	  ���           	 � ?  �  �  K         ����  t w          FJ� �       �   K   �   ��  �     	  ���           	 � �����  �  K         ����  ` c          Z\� �       �	  zX  >�   ��  �     
  ���           
 � >  �  �  W         ����  l n          `b� �       �	  �Y  "�   ��  �     
  ���           
 � ?  �  �  W         ����  { ~          fh� �       �	  �Z  �   ��  �     
  ���           
 � �����  �  W         ����  g h          ��� � t     �  �i  �   ��  �       ���            H  �  �  c         ����  s u          ��� � u     �  �j  �   ��  �       ���            I  �  �  c         ����  � �          ��� � v     �  *l  �   ��  �       ���            �����  �  c         ����  m o          ��� � ~     '  8|  �N   ��  �       ���            H  �  �  o         ����  z |          ��� �      V  �}   a   ��  �       ���            I  �  �  o         ����  � �          ��� � �     �    hs   ��  �       ���            �����  �  o         ����  p r          ��� � �     9  `�  @�   ��  �       ��0            R  �  �  �         ����  } �          ��� � �     p  �  ��   ��  �       ��0            S  �  �  �         ����  � �          ��� � �     �  l�  �   ��  �       ��0            �����  �  �         ����  x z          �� �     �  �  Һ	   ��  �       ��I            (R  �  �  �         ����  � �           �     '  ��  n�	   ��  �       ��I            'S  �  �  �         ����  � �          
�     f  V�  
�	   ��  �       ��I            &�����  �  �         ����  ~           5-2&�     H  B�   �   ��  �       ��J            5\  �  �  �         ����  � �          =58,�     �  �  @�   ��  �       ��J            4]  �  �  �         ����  � �          E=>2�     �  ��  `   ��  �       ��J            3�����  �  �         ����  U W          (� ~       E  p:  �   ��  ;       ��~            � 4  �  �  >         ����  ` a           .� �       [  `;  `   ��  ;       ��~            � 5  �  �  >         ����  m n          &4� �       q  P<  �   ��  ;       ��~            � �����  �  >         ����  [ ]          :G� �       @  �H   �   ��  <     	  ���           	 � >  �  �  J         ����  f h          @M� �       [  �I  ��   ��  <     	  ���           	 � ?  �  �  J         ����  t w          FS� �       v  �J  �   ��  <     	  ���           	 � �����  �  J         ����  ` c          Ze� �       �	  X  ��   ��  =     
  ���           
 � >  �  �  V         ����  l n          `k� �       �	  BY  ��   ��  =     
  ���           
 � ?  �  �  V         ����  { ~          fq� �       �	  nZ  ��   ��  =     
  ���           
 � �����  �  V         ����  g h          ��� � t     �  2i  X�   ��  >       ���            H  �  �  b         ����  s u          ��� � u     �  |j  ��   ��  >       ���            I  �  �  b         ����  � �          ��� � v     �  �k  H   ��  >       ���            �����  �  b         ����  m o          ��� � ~       �{  �I   ��  ?       ���            H  �  �  n         ����  z |          ��� �      I  <}  \   ��  ?       ���            I  �  �  n         ����  � �          ��� � �     x  �~  Tn   ��  ?       ���            �����  �  n         ����  p r          ��� � �     +  ��  ��   ��  @       ��6            R  �  �  �         ����  } �          ��� � �     b  ��  �   ��  @       ��6            S  �  �  �         ����  � �          ��� � �     �  �  p
   ��  @       ��6            �����  �  �         ����  x z          � �     �  ��  ��	   ��  A       ��U            (R  �  �  �         ����  � �          	�       N�  ��	   ��  A       ��U            'S  �  �  �         ����  � �          
�     W  �  .�	   ��  A       ��U            &�����  �  �         ����  ~           562&�     8  ޼  ��   ��  B       ��V            5\  �  �  �         ����  � �          =>8,�     �  ��   �   ��  B       ��V            4]  �  �  �         ����  � �          EF>2�     �  b�      ��  B       ��V            3�����  �  �         ����  U W          � ~       �  xA  8M   ��  �       ���            � 4  �  �  @         ����  ` a           "� �       �  hB  �U   ��  �       ���            � 5  �  �  @         ����  m n          &(� �         XC  ^   ��  �       ���            � �����  �  @         ����  Y [          :;� �       �  �O  P   ��  �     	  ���           	 � >  �  �  L         ����  c f          @A� �         �P  �%   ��  �     	  ���           	 � ?  �  �  L         ����  q t          FG� �       *  �Q  h0   ��  �     	  ���           	 � �����  �  L         ����  ` c          ZY� �       v
  _  J   ��  �     
  ���           
 � >  �  �  X         ����  l n          `_� �       �
  J`  .#   ��  �     
  ���           
 � ?  �  �  X         ����  { ~          fe� �       �
  va  0   ��  �     
  ���           
 � �����  �  X         ����  g h          ��� � t     z  :p  �B   ��  �       ���            H  �  �  d         ����  s u          ��� � u     �  �q  0R   ��  �       ���            I  �  �  d         ����  � �          ��� � v     �  �r  �a   ��  �       ���            �����  �  d         ����  m o          ��� � ~       ܂  ,�   ��  �       ���            H  �  �  p         ����  z |          ��� �      3  D�  t�   ��  �       ���            I  �  �  p         ����  � �          ��� � �     b  ��  ��   ��  �       ���            �����  �  p         ����  p r          ��� � �     '  �  8B   ��  �       ��;            R  �  �  �         ����  } �          ��� � �     ^  ��  �W   ��  �       ��;            S  �  �  �         ����  � �          ��� � �     �  �  �l   ��  �       ��;            �����  �  �         ����  x z          �� �     �  ��  n
   ��  �       ��a            (R  �  �  �         ����  � �          ��     &  V�  
7
   ��  �       ��a            'S  �  �  �         ����  � �          
�     e  ��  �O
   ��  �       ��a            &�����  �  �         ����  ~           5*2&�     X  ��  `>   ��  �       ��b            5\  �  �  �         ����  � �          =28,�     �  ��  �Z   ��  �       ��b            4]  �  �  �         ����  � �          E:>2�     �  j�  �v   ��  �       ��b            3�����  �  �         ����  Y [          3� ~       �  �?  (?   ��         ���            � 4  �  �  B         ����  c f           9� �       �  �@  �G   ��         ���            � 5  �  �  B         ����  q t          &?� �       �  �A  P   ��         ���            � �����  �  B         ����  _ `          :R� �       �  �M  �   ��         ���           	 � >  �  �  N         ����  k l          @X� �       �  O  <   ��         ���           	 � ?  �  �  N         ����  z {          F^� �         P  �    ��         ���           	 � �����  �  N         ����  c e          Zp� �       J
  �]     ��  	     	  ���           
 � >  �  �  Z         ����  n q          `v� �       k
  �^  �   ��  	     	  ���           
 � ?  �  �  Z         ����  ~ �          f|� �       �
  �_  �   ��  	     	  ���           
 � �����  �  Z         ����  h j          ��� � t     J  �n  �/   ��  
     
  ���            H  �  �  f         ����  u w          ��� � u     r  �o  p?   ��  
     
  ���            I  �  �  f         ����  � �          ��� � v     �  >q  �N   ��  
     
  ���            �����  �  f         ����  o p          ��� � ~     �  L�  ܐ   ��         ���            H  �  �  r         ����  | }          ��� �      �  ��  $�   ��         ���            I  �  �  r         ����  � �          ��� � �     .  �  l�   ��         ���            �����  �  r         ����  t v          ��� � �     �  t�  X,   ��         ��@            R  �  �  �         ����  � �          ��� � �     &  ��  �A   ��         ��@            S  �  �  �         ����  � �          ��� � �     ]  ��   W   ��         ��@            �����  �  �         ����  | ~          � �     �  "�  �
   ��         ��m            (R  �  �            ����  � �          �     �  Ƭ  �
   ��         ��m            'S  �  �            ����  � �          
�     )  j�  68
   ��         ��m            &�����  �            ����   �          5A2&�       V�  `%   ��         ��n            5\  �  �           ����  � �          =I8,�     `  �  �A   ��         ��n            4]  �  �           ����  � �          EQ>2�     �  ��  �]   ��         ��n            3�����  �           ����  W Y           � ~       �  X>  1   ��  m       ���            � 4  �  �  A         ����  a c           &� �       �  H?  �9   ��  m       ���            � 5  �  �  A         ����  n q          &,� �       �  8@  �A   ��  m       ���            � �����  �  A         ����  ] _          :?� �       �  hL  �   ��  n     	  ���           	 � >  �  �  M         ����  h k          @E� �       �  vM  �   ��  n     	  ���           	 � ?  �  �  M         ����  w z          FK� �       �  �N  (   ��  n     	  ���           	 � �����  �  M         ����  c e          Z]� �       
  �[  ��   ��  o     
  ���           
 � >  �  �  Y         ����  n q          `c� �       ?
  *]  �    ��  o     
  ���           
 � ?  �  �  Y         ����  ~ �          fi� �       `
  V^  �   ��  o     
  ���           
 � �����  �  Y         ����  h j          ��� � t       m  8   ��  p       ���            H  �  �  e         ����  u w          ��� � u     B  dn  �,   ��  p       ���            I  �  �  e         ����  � �          ��� � v     j  �o  (<   ��  p       ���            �����  �  e         ����  m o          ��� � ~     �  �  �|   ��  q       ���            H  �  �  q         ����  z |          ��� �      �  $�  Ԏ   ��  q       ���            I  �  �  q         ����  � �          ��� � �     �  ��  �   ��  q       ���            �����  �  q         ����  r t          ��� � �     �  �  x   ��  r       ��E            R  �  �  �         ����  � �          ��� � �     �  j�  �+   ��  r       ��E            S  �  �  �         ����  � �          ��� � �     %  �   A   ��  r       ��E            �����  �  �         ����  z |          �� �     o  ��  ��	   ��  s       ��y            (R  �  �           ����  � �          �     �  6�  *
   ��  s       ��y            'S  �  �           ����  � �          
�     �  ڬ  � 
   ��  s       ��y            &�����  �           ����   �          5.2&�     �  ��  `   ��  t       ��z            5\  �  �           ����  � �          =68,�        ��  �(   ��  t       ��z            4]  �  �           ����  � �          E>>2�     h  J�  �D   ��  t       ��z            3�����  �           ����    U W          � � l~       {  �<  #   ��         ��^            � 4  �  �  
         ����    ` a          � � s�       �  �=  x+   ��         ��^            � 5  �  �  
         ����    m n          � � z�       �  �>  �3   ��         ��^            � �����  �  
         ����    [ ]          � � ��       |  �J  p�   ��  �     	  ��_           	 � >  �  �           ����    f h          � � ��       �  �K  ��   ��  �     	  ��_           	 � ?  �  �           ����    t w          � � ��       �  �L  �   ��  �     	  ��_           	 � �����  �           ����    _ `          �  ��       �	  nZ  ��   ��  �     
  ��`           
 � >  �  �           ����    k l          � ��       
  �[  ��   ��  �     
  ��`           
 � ?  �  �           ����    z {          � 
��       4
  �\  ��   ��  �     
  ��`           
 � �����  �           ����    e g          � &�� t     �  �k  x
   ��  �       ��a            H  �  �           ����    q s          � ,�� u       �l  �   ��  �       ��a            I  �  �           ����    � �          � 2�� v     :  n  h)   ��  �       ��a            �����  �           ����    j m          � E� ~     h  ,~  <h   ��  �       ��b            H  �  �           ����    w z          � K"�      �  �  �z   ��  �       ��b            I  �  �           ����    � �          � Q*� �     �  ��  ̌   ��  �       ��b            �����  �           ����    p r          	cI� �       T�  �    ��  �       ��c            R  �  �           ����    } �          iQ� �     �  ړ  �   ��  �       ��c            S  �  �           ����    � �          oY� �     �  `�  @+   ��  �       ��c            �����  �           ����    x z          0�x �     3  �  �	   ��  �       ��?            (R  �  �  �         ����    � �          6���     r  ��  ��	   ��  �       ��?            'S  �  �  �         ����    � �          <��
�     �  J�  V	
   ��  �       ��?            &�����  �  �         ����    | ~          P��&�     �  6�  `�   ��  �       ��@            5\  �  �  �         ����    � �          V��,�     �  ��  �   ��  �       ��@            4]  �  �  �         ����    � �          \��2�     (  ��  �+   ��  �       ��@            3�����  �  �         ����   S U          � � `~       N  �:  t   ��  �       ��k            � 4  �  �           ����   ] `          � � g�       d  �;  �   ��  �       ��k            � 5  �  �           ����   j m          � � n�       z  �<  T"   ��  �       ��k            � �����  �           ����   Y [          � � ��       J  �H  ��   ��  �     	  ��l           	 � >  �  �           ����   c f          � � ��       e  �I  t�   ��  �     	  ��l           	 � ?  �  �           ����   q t          � � ��       �   K   �   ��  �     	  ��l           	 � �����  �           ����   _ `          �  ��       �	  zX  >�   ��  �     
  ��m           
 � >  �  �           ����   k l          � ��       �	  �Y  "�   ��  �     
  ��m           
 � ?  �  �           ����   z {          � 
��       �	  �Z  �   ��  �     
  ��m           
 � �����  �           ����   c e          � &�� t     �  �i  �   ��  �       ��n            H  �  �           ����   n q          � ,�� u     �  �j  �   ��  �       ��n            I  �  �           ����   ~ �          � 2�� v     �  *l  �   ��  �       ��n            �����  �           ����   h j          � E� ~     '  8|  �N   ��  �       ��o            H  �  �           ����   u w          � K�      V  �}   a   ��  �       ��o            I  �  �           ����   � �          � Q� �     �    hs   ��  �       ��o            �����  �           ����   o p          	c=� �     9  `�  @�   ��  �       ��p            R  �  �           ����   | }          iE� �     p  �  ��   ��  �       ��p            S  �  �           ����   � �          oM� �     �  l�  �   ��  �       ��p            �����  �           ����   v x          0�l �     �  �  Һ	   ��  �       ��K            (R  �  �  �         ����   � �          6�t�     '  ��  n�	   ��  �       ��K            'S  �  �  �         ����   � �          <�|
�     f  V�  
�	   ��  �       ��K            &�����  �  �         ����   | ~          P��&�     H  B�   �   ��  �       ��L            5\  �  �  �         ����   � �          V��,�     �  �  @�   ��  �       ��L            4]  �  �  �         ����   � �          \��2�     �  ��  `   ��  �       ��L            3�����  �  �         ����   S U          � � h~       E  p:  �   ��  L       ��x            � 4  �  �  $         ����   ] `          � � o�       [  `;  `   ��  L       ��x            � 5  �  �  $         ����   j m          � � v�       q  P<  �   ��  L       ��x            � �����  �  $         ����   Y [          � � ��       @  �H   �   ��  M     	  ��y           	 � >  �  �  %         ����   c f          � � ��       [  �I  ��   ��  M     	  ��y           	 � ?  �  �  %         ����   q t          � � ��       v  �J  �   ��  M     	  ��y           	 � �����  �  %         ����   _ `          �  ��       �	  X  ��   ��  N     
  ��z           
 � >  �  �  &         ����   k l          � ��       �	  BY  ��   ��  N     
  ��z           
 � ?  �  �  &         ����   z {          � 
��       �	  nZ  ��   ��  N     
  ��z           
 � �����  �  &         ����   c e          � &�� t     �  2i  X�   ��  O       ��{            H  �  �  '         ����   n q          � ,�� u     �  |j  ��   ��  O       ��{            I  �  �  '         ����   ~ �          � 2�� v     �  �k  H   ��  O       ��{            �����  �  '         ����   h j          � E� ~       �{  �I   ��  P       ��|            H  �  �  (         ����   u w          � K�      I  <}  \   ��  P       ��|            I  �  �  (         ����   � �          � Q&� �     x  �~  Tn   ��  P       ��|            �����  �  (         ����   o p          	cE� �     +  ��  ��   ��  Q       ��}            R  �  �  )         ����   | }          iM� �     b  ��  �   ��  Q       ��}            S  �  �  )         ����   � �          oU� �     �  �  p
   ��  Q       ��}            �����  �  )         ����   v x          0�t �     �  ��  ��	   ��  R       ��W            (R  �  �  �         ����   � �          6�|�       N�  ��	   ��  R       ��W            'S  �  �  �         ����   � �          <��
�     W  �  .�	   ��  R       ��W            &�����  �  �         ����   | ~          P��&�     8  ޼  ��   ��  S       ��X            5\  �  �  �         ����   � �          V��,�     �  ��   �   ��  S       ��X            4]  �  �  �         ����   � �          \��2�     �  b�      ��  S       ��X            3�����  �  �         ����   S U          � � \~       �  xA  8M   ��  �       ���            � 4  �  �  1         ����   ] `          � � c�       �  hB  �U   ��  �       ���            � 5  �  �  1         ����   j m          � � j�         XC  ^   ��  �       ���            � �����  �  1         ����   Y [          � � ��       �  �O  P   ��  �     	  ���           	 � >  �  �  2         ����   c f          � � ��         �P  �%   ��  �     	  ���           	 � ?  �  �  2         ����   q t          � � ��       *  �Q  h0   ��  �     	  ���           	 � �����  �  2         ����   _ `          �  ��       v
  _  J   ��  �     
  ���           
 � >  �  �  3         ����   k l          � ��       �
  J`  .#   ��  �     
  ���           
 � ?  �  �  3         ����   z {          � 
��       �
  va  0   ��  �     
  ���           
 � �����  �  3         ����   c e          � &�� t     z  :p  �B   ��  �       ���            H  �  �  4         ����   n q          � ,�� u     �  �q  0R   ��  �       ���            I  �  �  4         ����   ~ �          � 2�� v     �  �r  �a   ��  �       ���            �����  �  4         ����   h j          � E
� ~       ܂  ,�   ��  �       ���            H  �  �  5         ����   u w          � K�      3  D�  t�   ��  �       ���            I  �  �  5         ����   � �          � Q� �     b  ��  ��   ��  �       ���            �����  �  5         ����   o p          	c9� �     '  �  8B   ��  �       ���            R  �  �  6         ����   | }          iA� �     ^  ��  �W   ��  �       ���            S  �  �  6         ����   � �          oI� �     �  �  �l   ��  �       ���            �����  �  6         ����   v x          0�h �     �  ��  n
   ��  �       ��c            (R  �  �  �         ����   � �          6�p�     &  V�  
7
   ��  �       ��c            'S  �  �  �         ����   � �          <�x
�     e  ��  �O
   ��  �       ��c            &�����  �  �         ����   | ~          P��&�     X  ��  `>   ��  �       ��d            5\  �  �  �         ����   � �          V��,�     �  ��  �Z   ��  �       ��d            4]  �  �  �         ����   � �          \��2�     �  j�  �v   ��  �       ��d            3�����  �  �         ����   U W          � � t~       �  �?  (?   ��         ���            � 4  �  �  >         ����   ` a          � � {�       �  �@  �G   ��         ���            � 5  �  �  >         ����   m n          � � ��       �  �A  P   ��         ���            � �����  �  >         ����   [ ]          � � ��       �  �M  �   ��         ���           	 � >  �  �  ?         ����   f h          � � ��       �  O  <   ��         ���           	 � ?  �  �  ?         ����   t w          � � ��         P  �    ��         ���           	 � �����  �  ?         ����   _ `          �  ��       J
  �]     ��       	  ���           
 � >  �  �  @         ����   k l          � ��       k
  �^  �   ��       	  ���           
 � ?  �  �  @         ����   z {          � 
��       �
  �_  �   ��       	  ���           
 � �����  �  @         ����   e g          � &�� t     J  �n  �/   ��       
  ���            H  �  �  A         ����   q s          � ,�� u     r  �o  p?   ��       
  ���            I  �  �  A         ����   � �          � 2�� v     �  >q  �N   ��       
  ���            �����  �  A         ����   j m          � E"� ~     �  L�  ܐ   ��         ���            H  �  �  B         ����   w z          � K*�      �  ��  $�   ��         ���            I  �  �  B         ����   � �          � Q2� �     .  �  l�   ��         ���            �����  �  B         ����   p r          	cQ� �     �  t�  X,   ��         ���            R  �  �  C         ����   } �          iY� �     &  ��  �A   ��         ���            S  �  �  C         ����   � �          oa� �     ]  ��   W   ��         ���            �����  �  C         ����   x z          0�� �     �  "�  �
   ��         ��o            (R  �  �           ����   � �          6���     �  Ƭ  �
   ��         ��o            'S  �  �           ����   � �          <��
�     )  j�  68
   ��         ��o            &�����  �           ����   | ~          P��&�       V�  `%   ��         ��p            5\  �  �           ����   � �          V��,�     `  �  �A   ��         ��p            4]  �  �           ����   � �          \��2�     �  ��  �]   ��         ��p            3�����  �           ����   S U          � � d~       �  X>  1   ��  ~       ���            � 4  �  �  K         ����   ] `          � � k�       �  H?  �9   ��  ~       ���            � 5  �  �  K         ����   j m          � � r�       �  8@  �A   ��  ~       ���            � �����  �  K         ����   Y [          � � ��       �  hL  �   ��       	  ���           	 � >  �  �  L         ����   c f          � � ��       �  vM  �   ��       	  ���           	 � ?  �  �  L         ����   q t          � � ��       �  �N  (   ��       	  ���           	 � �����  �  L         ����   _ `          �  ��       
  �[  ��   ��  �     
  ���           
 � >  �  �  M         ����   k l          � ��       ?
  *]  �    ��  �     
  ���           
 � ?  �  �  M         ����   z {          � 
��       `
  V^  �   ��  �     
  ���           
 � �����  �  M         ����   c e          � &�� t       m  8   ��  �       ���            H  �  �  N         ����   n q          � ,�� u     B  dn  �,   ��  �       ���            I  �  �  N         ����   ~ �          � 2�� v     j  �o  (<   ��  �       ���            �����  �  N         ����   h j          � E� ~     �  �  �|   ��  �       ���            H  �  �  O         ����   u w          � K�      �  $�  Ԏ   ��  �       ���            I  �  �  O         ����   � �          � Q"� �     �  ��  �   ��  �       ���            �����  �  O         ����   o p          	cA� �     �  �  x   ��  �       ���            R  �  �  P         ����   | }          iI� �     �  j�  �+   ��  �       ���            S  �  �  P         ����   � �          oQ� �     %  �   A   ��  �       ���            �����  �  P         ����   v x          0�p �     o  ��  ��	   ��  �       ��{            (R  �  �           ����   � �          6�x�     �  6�  *
   ��  �       ��{            'S  �  �           ����   � �          <��
�     �  ڬ  � 
   ��  �       ��{            &�����  �           ����   | ~          P��&�     �  ��  `   ��  �       ��|            5\  �  �           ����   � �          V��,�        ��  �(   ��  �       ��|            4]  �  �           ����   � �          \��2�     h  J�  �D   ��  �       ��|            3�����  �           ����   U W          � � p~         C  H[   ��  �     �   �            � 4  �  �  X         ����   ` a          � � w�       !  �C  �c   ��  �     �   �            � 5  �  �  X         ����   m n          � � ~�       7  �D  (l   ��  �     �   �            � �����  �  X         ����   [ ]          � � ��         Q  �*   ��  �     �   �           	 � >  �  �  Y         ����   f h          � � ��       7  &R  |5   ��  �     �   �           	 � ?  �  �  Y         ����   t w          � � ��       R  4S  @   ��  �     �   �           	 � �����  �  Y         ����   _ `          �  ��       �
  �`  z'   ��  �     �   �           
 � >  �  �  Z         ����   k l          � ��       �
  �a  ^4   ��  �     �   �           
 � ?  �  �  Z         ����   z {          � 
��       �
  c  BA   ��  �     �   �           
 � �����  �  Z         ����   e g          � &�� t     �  �q  xU   ��  �     �   �            H  �  �  [         ����   q s          � ,�� u     �  s  �d   ��  �     �   �            I  �  �  [         ����   � �          � 2�� v     �  ^t  ht   ��  �     �   �            �����  �  [         ����   j m          � E� ~     8  l�  |�   ��  �     �   �            H  �  �  \         ����   w z          � K&�      g  ԅ  ��   ��  �     �   �            I  �  �  \         ����   � �          � Q.� �     �  <�  �   ��  �     �   �            �����  �  \         ����   p r          	cM� �     _  ��  X   ��  �     �   �            R  �  �  ]         ����   } �          iU� �     �  �  lm   ��  �     �   �            S  �  �  ]         ����   � �          o]� �     �  ��  ��   ��  �     �   �            �����  �  ]         ����   x z          0�| �     #  B�  �5
   ��  �     �   �            (R  �  �           ����   � �          6���     b  �  zN
   ��  �     �   �            'S  �  �           ����   � �          <��
�     �  ��  g
   ��  �     �   �            &�����  �           ����   | ~          P��&�     �  v�  `W   ��  �     �   �            5\  �  �           ����   � �          V��,�     �  8�  �s   ��  �     �   �            4]  �  �           ����   � �          \��2�     (   ��  ��   ��  �     �   �            3�����  �        